# 
# LEF OUT 
# User Name : islam 
# Date : Mon May  9 14:20:45 2022
# 
VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 10000 ;
END UNITS
MANUFACTURINGGRID 0.0005 ;

LAYER active
  TYPE MASTERSLICE ;
  MASK 3 ;
END active

LAYER nwell
  TYPE MASTERSLICE ;
  MASK 3 ;
END nwell

LAYER m1text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m1text

LAYER m2text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m2text

LAYER m3text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m3text

LAYER m4text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m4text

LAYER m5text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m5text

LAYER m6text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m6text

LAYER m7text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m7text

LAYER m8text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m8text

LAYER m9text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m9text

LAYER m10text
  TYPE MASTERSLICE ;
  MASK 3 ;
END m10text

LAYER pimplant
  TYPE MASTERSLICE ;
  MASK 3 ;
END pimplant

LAYER nimplant
  TYPE MASTERSLICE ;
  MASK 3 ;
END nimplant

LAYER outline
  TYPE MASTERSLICE ;
  MASK 3 ;
END outline

LAYER metal1
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.14 ;
  WIDTH 0.065 ;
  AREA 0.01 ;
  SPACING   0.065 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.065 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 85 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 60 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal1

LAYER via1
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.075 ;
  WIDTH 0.065 ;
END via1

LAYER metal2
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION VERTICAL ;
  PITCH 0.19 ;
  WIDTH 0.07 ;
  AREA 0.01 ;
  SPACING   0.07 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.07 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal2

LAYER via2
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.38 ;
  WIDTH 0.07 ;
  AREA 0.01 ;
  SPACING   0.07 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.07 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal3

LAYER via3
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.085 ;
  WIDTH 0.07 ;
END via3

LAYER metal4
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION VERTICAL ;
  PITCH 0.38 ;
  WIDTH 0.14 ;
  OFFSET 0.19 ;
  AREA 0.01 ;
  SPACING   0.14 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.14 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal4

LAYER via4
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
END via4

LAYER metal5
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION HORIZONTAL ;
  PITCH 0.76 ;
  WIDTH 0.14 ;
  AREA 0.01 ;
  SPACING   0.14 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.14 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal5

LAYER via5
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
END via5

LAYER metal6
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION VERTICAL ;
  PITCH 0.76 ;
  WIDTH 0.14 ;
  OFFSET 0.38 ;
  AREA 0.01 ;
  SPACING   0.14 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.14 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal6

LAYER via6
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.16 ;
  WIDTH 0.14 ;
END via6

LAYER metal7
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION HORIZONTAL ;
  PITCH 1.52 ;
  WIDTH 0.4 ;
  AREA 0.01 ;
  SPACING   0.4 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.4 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal7

LAYER via7
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
END via7

LAYER metal8
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION VERTICAL ;
  PITCH 1.52 ;
  WIDTH 0.4 ;
  OFFSET 0.76 ;
  AREA 0.01 ;
  SPACING   0.4 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.4 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal8

LAYER via8
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.44 ;
  WIDTH 0.4 ;
END via8

LAYER metal9
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION HORIZONTAL ;
  PITCH 3.04 ;
  WIDTH 0.8 ;
  AREA 0.01 ;
  SPACING   0.8 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.8 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 60 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal9

LAYER via9
  TYPE CUT ;
  MASK 3 ;
  SPACING 0.88 ;
  WIDTH 0.8 ;
END via9

LAYER metal10
  TYPE ROUTING ;
  MASK 3 ;
  DIRECTION VERTICAL ;
  PITCH 3.04 ;
  WIDTH 0.8 ;
  OFFSET 1.52 ;
  AREA 0.01 ;
  SPACING   0.8 SAMENET ;
  MAXWIDTH 5 ;
  MINWIDTH 0.8 ;
  MINENCLOSEDAREA 0.2 ;
  CAPMULTIPLIER 1 ;
  MINIMUMDENSITY 15 ;
  MAXIMUMDENSITY 100 ;
  DENSITYCHECKWINDOW 50 50 ;
  DENSITYCHECKSTEP 25 ;
  MINIMUMDENSITY 1 ;
  MAXIMUMDENSITY 60 ;
  DENSITYCHECKWINDOW 100.00000 100.00000 ;
  DENSITYCHECKSTEP 50 ;
END metal10

LAYER OverlapCheck
  TYPE OVERLAP ;
END OverlapCheck

VIA VIA12
  DEFAULT 
  RESISTANCE 5.7 ;
  LAYER metal1 ;
    RECT -0.032500 -0.067500 0.032500 0.067500 ;
  LAYER via1 ;
    RECT -0.032500 -0.032500 0.032500 0.032500 ;
  LAYER metal2 ;
    RECT -0.067500 -0.032500 0.067500 0.032500 ;
END VIA12

VIA VIA23
  DEFAULT 
  RESISTANCE 5 ;
  LAYER metal2 ;
    RECT -0.070000 -0.035000 0.070000 0.035000 ;
  LAYER via2 ;
    RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal3 ;
    RECT -0.035000 -0.070000 0.035000 0.070000 ;
END VIA23

VIA VIA34
  DEFAULT 
  RESISTANCE 5 ;
  LAYER metal3 ;
    RECT -0.035000 -0.070000 0.035000 0.070000 ;
  LAYER via3 ;
    RECT -0.035000 -0.035000 0.035000 0.035000 ;
  LAYER metal4 ;
    RECT -0.035000 -0.035000 0.035000 0.035000 ;
END VIA34

VIA VIA45
  DEFAULT 
  RESISTANCE 3 ;
  LAYER metal4 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
  LAYER via4 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
  LAYER metal5 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
END VIA45

VIA VIA56
  DEFAULT 
  RESISTANCE 3 ;
  LAYER metal5 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
  LAYER via5 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
  LAYER metal6 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
END VIA56

VIA VIA67
  DEFAULT 
  RESISTANCE 3 ;
  LAYER metal6 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
  LAYER via6 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
  LAYER metal7 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
END VIA67

VIA VIA78
  DEFAULT 
  RESISTANCE 1 ;
  LAYER metal7 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
  LAYER via7 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
  LAYER metal8 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
END VIA78

VIA VIA89
  DEFAULT 
  RESISTANCE 1 ;
  LAYER metal8 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
  LAYER via8 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
  LAYER metal9 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
END VIA89

VIA VIA910
  DEFAULT 
  RESISTANCE 0.5 ;
  LAYER metal9 ;
    RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER via9 ;
    RECT -0.400000 -0.400000 0.400000 0.400000 ;
  LAYER metal10 ;
    RECT -0.400000 -0.400000 0.400000 0.400000 ;
END VIA910

VIARULE VIA12 GENERATE
  DEFAULT 
  LAYER metal1 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER via1 ;
    RECT -0.032500 -0.032500 0.032500 0.032500 ;
    SPACING 0.14 BY 0.14 ;
    RESISTANCE 5.7 ;
END VIA12

VIARULE VIA23 GENERATE
  DEFAULT 
  LAYER metal2 ;
    ENCLOSURE 0.035 0 ;
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER via2 ;
    RECT -0.035000 -0.035000 0.035000 0.035000 ;
    SPACING 0.155 BY 0.155 ;
    RESISTANCE 5 ;
END VIA23

VIARULE VIA34 GENERATE
  DEFAULT 
  LAYER metal3 ;
    ENCLOSURE 0 0.035 ;
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER via3 ;
    RECT -0.035000 -0.035000 0.035000 0.035000 ;
    SPACING 0.155 BY 0.155 ;
    RESISTANCE 5 ;
END VIA34

VIARULE VIA45 GENERATE
  DEFAULT 
  LAYER metal4 ;
    ENCLOSURE 0 0 ;
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER via4 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
    SPACING 0.3 BY 0.3 ;
    RESISTANCE 3 ;
END VIA45

VIARULE VIA56 GENERATE
  DEFAULT 
  LAYER metal5 ;
    ENCLOSURE 0 0 ;
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER via5 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
    SPACING 0.3 BY 0.3 ;
    RESISTANCE 3 ;
END VIA56

VIARULE VIA67 GENERATE
  DEFAULT 
  LAYER metal6 ;
    ENCLOSURE 0 0 ;
  LAYER metal7 ;
    ENCLOSURE 0.13 0.13 ;
  LAYER via6 ;
    RECT -0.070000 -0.070000 0.070000 0.070000 ;
    SPACING 0.3 BY 0.3 ;
    RESISTANCE 3 ;
END VIA67

VIARULE VIA78 GENERATE
  DEFAULT 
  LAYER metal7 ;
    ENCLOSURE 0 0 ;
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER via7 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
    SPACING 0.84 BY 0.84 ;
    RESISTANCE 1 ;
END VIA78

VIARULE VIA89 GENERATE
  DEFAULT 
  LAYER metal8 ;
    ENCLOSURE 0 0 ;
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER via8 ;
    RECT -0.200000 -0.200000 0.200000 0.200000 ;
    SPACING 0.84 BY 0.84 ;
    RESISTANCE 1 ;
END VIA89

VIARULE VIA910 GENERATE
  DEFAULT 
  LAYER metal9 ;
    ENCLOSURE 0 0 ;
  LAYER metal10 ;
    ENCLOSURE 0 0 ;
  LAYER via9 ;
    RECT -0.400000 -0.400000 0.400000 0.400000 ;
    SPACING 1.68 BY 1.68 ;
    RESISTANCE 0.5 ;
END VIA910

SITE unit
  CLASS CORE ;
  SYMMETRY X Y ;
  SIZE 0.19 BY 1.4 ;
END unit

MACRO XNOR2_X1
  CLASS CORE ;
  FOREIGN XNOR2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185000 0.390000 0.720000 0.460000 ;
        RECT 0.650000 0.460000 0.720000 0.555000 ;
        RECT 0.185000 0.460000 0.320000 0.560000 ;
        RECT 0.650000 0.555000 0.810000 0.625000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0688 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.350000 0.840000 0.965000 0.910000 ;
        RECT 0.350000 0.910000 0.510000 0.980000 ;
        RECT 0.895000 0.525000 0.965000 0.840000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0763 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2782 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END B

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.980000 1.100000 1.050000 ;
        RECT 0.630000 1.050000 0.700000 1.250000 ;
        RECT 1.030000 0.365000 1.100000 0.980000 ;
        RECT 0.785000 0.295000 1.100000 0.365000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.112 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4342 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.050000 1.115000 0.120000 1.315000 ;
        RECT 0.430000 1.115000 0.500000 1.315000 ;
        RECT 1.000000 1.115000 1.070000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.395000 0.085000 0.530000 0.250000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.210000 1.145000 0.345000 1.215000 ;
      RECT 0.210000 0.740000 0.280000 1.145000 ;
      RECT 0.050000 0.670000 0.585000 0.740000 ;
      RECT 0.515000 0.525000 0.585000 0.670000 ;
      RECT 0.050000 0.150000 0.120000 0.670000 ;
      RECT 0.595000 0.160000 1.105000 0.230000 ;
  END
END XNOR2_X1

MACRO XNOR2_X2
  CLASS CORE ;
  FOREIGN XNOR2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.15675 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal2 ;
    ANTENNAGATEAREA 0.15675 LAYER metal3 ;
    ANTENNAGATEAREA 0.15675 LAYER metal4 ;
    ANTENNAGATEAREA 0.15675 LAYER metal5 ;
    ANTENNAGATEAREA 0.15675 LAYER metal6 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ;
    ANTENNAGATEAREA 0.15675 LAYER metal8 ;
    ANTENNAGATEAREA 0.15675 LAYER metal9 ;
    ANTENNAGATEAREA 0.15675 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.505000 0.560000 0.890000 0.630000 ;
        RECT 0.820000 0.630000 0.890000 0.770000 ;
        RECT 0.820000 0.770000 1.650000 0.840000 ;
        RECT 1.580000 0.525000 1.650000 0.770000 ;
    END
    ANTENNAGATEAREA 0.15675 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.112 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4342 LAYER metal1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal2 ;
    ANTENNAGATEAREA 0.15675 LAYER metal3 ;
    ANTENNAGATEAREA 0.15675 LAYER metal4 ;
    ANTENNAGATEAREA 0.15675 LAYER metal5 ;
    ANTENNAGATEAREA 0.15675 LAYER metal6 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ;
    ANTENNAGATEAREA 0.15675 LAYER metal8 ;
    ANTENNAGATEAREA 0.15675 LAYER metal9 ;
    ANTENNAGATEAREA 0.15675 LAYER metal10 ;
  END B

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.210000 0.905000 1.840000 0.975000 ;
        RECT 1.770000 0.430000 1.840000 0.905000 ;
        RECT 0.975000 0.360000 1.840000 0.430000 ;
        RECT 1.765000 0.190000 1.840000 0.360000 ;
    END
    ANTENNADIFFAREA 0.32165 ;
    ANTENNAPARTIALMETALAREA 0.22065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8346 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.900000 1.485000 ;
        RECT 1.540000 1.240000 1.675000 1.315000 ;
        RECT 0.050000 1.065000 0.120000 1.315000 ;
        RECT 0.425000 1.065000 0.495000 1.315000 ;
        RECT 0.805000 1.065000 0.875000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.900000 0.085000 ;
        RECT 0.050000 0.085000 0.120000 0.325000 ;
        RECT 0.395000 0.085000 0.530000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.245000 0.725000 0.720000 0.795000 ;
      RECT 0.245000 0.460000 0.315000 0.725000 ;
      RECT 0.245000 0.390000 0.910000 0.460000 ;
      RECT 0.210000 0.225000 1.675000 0.295000 ;
      RECT 0.975000 1.095000 1.865000 1.165000 ;
  END
END XNOR2_X2

MACRO XOR2_X1
  CLASS CORE ;
  FOREIGN XOR2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.175000 0.665000 0.245000 0.730000 ;
        RECT 0.175000 0.730000 0.700000 0.800000 ;
        RECT 0.630000 0.660000 0.700000 0.730000 ;
        RECT 0.630000 0.525000 0.755000 0.660000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.063075 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2392 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.305000 0.875000 0.890000 0.945000 ;
        RECT 0.820000 0.660000 0.890000 0.875000 ;
        RECT 0.820000 0.525000 0.945000 0.660000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.072875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2756 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END B

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.775000 1.040000 1.080000 1.110000 ;
        RECT 1.010000 0.420000 1.080000 1.040000 ;
        RECT 0.620000 0.350000 1.080000 0.420000 ;
        RECT 0.620000 0.150000 0.690000 0.350000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.11095 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4303 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.420000 1.150000 0.490000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.285000 ;
        RECT 0.420000 0.085000 0.490000 0.285000 ;
        RECT 0.990000 0.085000 1.060000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.040000 0.595000 0.110000 1.250000 ;
      RECT 0.040000 0.525000 0.565000 0.595000 ;
      RECT 0.495000 0.595000 0.565000 0.660000 ;
      RECT 0.225000 0.150000 0.295000 0.525000 ;
      RECT 0.585000 1.175000 1.095000 1.245000 ;
  END
END XOR2_X1

MACRO XOR2_X2
  CLASS CORE ;
  FOREIGN XOR2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.285000 0.820000 0.355000 ;
        RECT 0.745000 0.355000 0.820000 0.395000 ;
        RECT 0.060000 0.355000 0.165000 0.700000 ;
        RECT 0.745000 0.395000 1.325000 0.465000 ;
        RECT 0.745000 0.465000 0.820000 0.660000 ;
        RECT 1.255000 0.465000 1.325000 0.660000 ;
    END
    ANTENNAGATEAREA 0.15675 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1613 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5668 LAYER metal1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal2 ;
    ANTENNAGATEAREA 0.15675 LAYER metal3 ;
    ANTENNAGATEAREA 0.15675 LAYER metal4 ;
    ANTENNAGATEAREA 0.15675 LAYER metal5 ;
    ANTENNAGATEAREA 0.15675 LAYER metal6 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ;
    ANTENNAGATEAREA 0.15675 LAYER metal8 ;
    ANTENNAGATEAREA 0.15675 LAYER metal9 ;
    ANTENNAGATEAREA 0.15675 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.365000 0.560000 0.500000 0.770000 ;
        RECT 0.365000 0.770000 1.125000 0.840000 ;
        RECT 0.990000 0.560000 1.125000 0.770000 ;
    END
    ANTENNAGATEAREA 0.15675 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1099 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER metal1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal2 ;
    ANTENNAGATEAREA 0.15675 LAYER metal3 ;
    ANTENNAGATEAREA 0.15675 LAYER metal4 ;
    ANTENNAGATEAREA 0.15675 LAYER metal5 ;
    ANTENNAGATEAREA 0.15675 LAYER metal6 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ;
    ANTENNAGATEAREA 0.15675 LAYER metal8 ;
    ANTENNAGATEAREA 0.15675 LAYER metal9 ;
    ANTENNAGATEAREA 0.15675 LAYER metal10 ;
  END B

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.800000 0.905000 1.465000 0.975000 ;
        RECT 1.390000 0.330000 1.465000 0.905000 ;
        RECT 0.885000 0.260000 1.465000 0.330000 ;
        RECT 0.885000 0.220000 0.955000 0.260000 ;
        RECT 0.610000 0.150000 0.955000 0.220000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.157225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5902 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.445000 1.205000 0.515000 1.315000 ;
        RECT 1.585000 1.205000 1.655000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.070000 0.085000 0.140000 0.210000 ;
        RECT 0.445000 0.085000 0.515000 0.195000 ;
        RECT 1.025000 0.085000 1.095000 0.195000 ;
        RECT 1.585000 0.085000 1.655000 0.335000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.610000 1.175000 1.500000 1.245000 ;
      RECT 0.040000 1.040000 1.600000 1.110000 ;
      RECT 1.530000 0.525000 1.600000 1.040000 ;
      RECT 0.230000 0.495000 0.300000 1.040000 ;
      RECT 0.230000 0.425000 0.645000 0.495000 ;
      RECT 0.575000 0.495000 0.645000 0.660000 ;
  END
END XOR2_X2

MACRO TAP
  CLASS CORE ;
  FOREIGN TAP 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.380000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.380000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
    END
  END VSS
END TAP

MACRO OAI22_X4
  CLASS CORE ;
  FOREIGN OAI22_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.910000 0.560000 2.045000 0.725000 ;
        RECT 1.910000 0.725000 2.805000 0.795000 ;
        RECT 2.670000 0.560000 2.805000 0.725000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1072 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3367 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.645000 0.425000 3.035000 0.495000 ;
        RECT 1.645000 0.495000 1.715000 0.660000 ;
        RECT 2.320000 0.495000 2.390000 0.660000 ;
        RECT 2.910000 0.495000 3.035000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.146025 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5187 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.560000 0.520000 0.725000 ;
        RECT 0.385000 0.725000 1.280000 0.795000 ;
        RECT 1.145000 0.560000 1.280000 0.725000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1072 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3367 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.150000 0.425000 1.520000 0.495000 ;
        RECT 0.150000 0.495000 0.220000 0.660000 ;
        RECT 0.795000 0.495000 0.865000 0.660000 ;
        RECT 1.390000 0.495000 1.520000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.14565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5135 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.865000 3.170000 0.935000 ;
        RECT 0.425000 0.935000 0.495000 1.210000 ;
        RECT 1.175000 0.935000 1.245000 1.210000 ;
        RECT 1.935000 0.935000 2.005000 1.210000 ;
        RECT 2.695000 0.935000 2.765000 1.210000 ;
        RECT 3.100000 0.360000 3.170000 0.865000 ;
        RECT 1.720000 0.290000 3.170000 0.360000 ;
    END
    ANTENNADIFFAREA 0.5852 ;
    ANTENNAPARTIALMETALAREA 0.406 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5262 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.230000 1.485000 ;
        RECT 0.040000 1.040000 0.110000 1.315000 ;
        RECT 0.795000 1.040000 0.865000 1.315000 ;
        RECT 1.555000 1.040000 1.625000 1.315000 ;
        RECT 2.315000 1.040000 2.385000 1.315000 ;
        RECT 3.075000 1.040000 3.145000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.230000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.195000 ;
        RECT 0.605000 0.085000 0.675000 0.195000 ;
        RECT 0.985000 0.085000 1.055000 0.195000 ;
        RECT 1.365000 0.085000 1.435000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.260000 1.595000 0.330000 ;
      RECT 1.525000 0.220000 1.595000 0.260000 ;
      RECT 0.045000 0.185000 0.115000 0.260000 ;
      RECT 1.525000 0.150000 3.180000 0.220000 ;
  END
END OAI22_X4

MACRO OAI33_X1
  CLASS CORE ;
  FOREIGN OAI33_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145000 0.525000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.365000 1.260000 0.435000 ;
        RECT 0.630000 0.435000 0.700000 1.000000 ;
        RECT 1.190000 0.150000 1.260000 0.365000 ;
    END
    ANTENNADIFFAREA 0.189875 ;
    ANTENNAPARTIALMETALAREA 0.0987 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3848 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.055000 0.975000 0.125000 1.315000 ;
        RECT 1.190000 0.975000 1.260000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.335000 ;
        RECT 0.400000 0.085000 0.535000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215000 0.225000 1.105000 0.295000 ;
  END
END OAI33_X1

MACRO OR2_X1
  CLASS CORE ;
  FOREIGN OR2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.610000 0.150000 0.700000 1.240000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0981 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3068 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.415000 0.965000 0.485000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.285000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.900000 0.115000 1.240000 ;
      RECT 0.045000 0.830000 0.540000 0.900000 ;
      RECT 0.470000 0.420000 0.540000 0.830000 ;
      RECT 0.235000 0.350000 0.540000 0.420000 ;
      RECT 0.235000 0.150000 0.305000 0.350000 ;
  END
END OR2_X1

MACRO OR2_X2
  CLASS CORE ;
  FOREIGN OR2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615000 0.150000 0.700000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.415000 1.040000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.975000 0.115000 1.250000 ;
      RECT 0.045000 0.905000 0.545000 0.975000 ;
      RECT 0.475000 0.425000 0.545000 0.905000 ;
      RECT 0.235000 0.355000 0.545000 0.425000 ;
      RECT 0.235000 0.150000 0.305000 0.355000 ;
  END
END OR2_X2

MACRO OR2_X4
  CLASS CORE ;
  FOREIGN OR2_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.150000 0.765000 ;
        RECT 0.060000 0.765000 0.760000 0.835000 ;
        RECT 0.690000 0.525000 0.760000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0874 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.150000 1.075000 0.560000 ;
        RECT 0.995000 0.560000 1.435000 0.700000 ;
        RECT 0.995000 0.700000 1.065000 1.095000 ;
        RECT 1.365000 0.700000 1.435000 1.095000 ;
        RECT 1.365000 0.150000 1.435000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1784 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5694 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.040000 1.035000 0.110000 1.315000 ;
        RECT 0.795000 1.035000 0.865000 1.315000 ;
        RECT 1.175000 1.035000 1.245000 1.315000 ;
        RECT 1.555000 1.035000 1.625000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.285000 ;
        RECT 1.175000 0.085000 1.245000 0.425000 ;
        RECT 1.555000 0.085000 1.625000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.425000 0.970000 0.495000 1.250000 ;
      RECT 0.425000 0.900000 0.925000 0.970000 ;
      RECT 0.855000 0.425000 0.925000 0.900000 ;
      RECT 0.235000 0.355000 0.925000 0.425000 ;
      RECT 0.235000 0.150000 0.305000 0.355000 ;
      RECT 0.605000 0.150000 0.675000 0.355000 ;
  END
END OR2_X4

MACRO OR3_X1
  CLASS CORE ;
  FOREIGN OR3_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.570000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.800000 0.150000 0.890000 1.240000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0981 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3068 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.605000 0.965000 0.675000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.900000 0.115000 1.240000 ;
      RECT 0.045000 0.830000 0.730000 0.900000 ;
      RECT 0.660000 0.420000 0.730000 0.830000 ;
      RECT 0.045000 0.350000 0.730000 0.420000 ;
      RECT 0.045000 0.150000 0.115000 0.350000 ;
      RECT 0.415000 0.150000 0.485000 0.350000 ;
  END
END OR3_X1

MACRO OR3_X2
  CLASS CORE ;
  FOREIGN OR3_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.570000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805000 0.150000 0.890000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.605000 0.975000 0.675000 1.315000 ;
        RECT 0.985000 0.975000 1.055000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
        RECT 0.985000 0.085000 1.055000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.910000 0.115000 1.250000 ;
      RECT 0.045000 0.840000 0.730000 0.910000 ;
      RECT 0.660000 0.460000 0.730000 0.840000 ;
      RECT 0.045000 0.390000 0.730000 0.460000 ;
      RECT 0.045000 0.150000 0.115000 0.390000 ;
      RECT 0.415000 0.150000 0.485000 0.390000 ;
  END
END OR3_X2

MACRO OR3_X4
  CLASS CORE ;
  FOREIGN OR3_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.610000 0.560000 0.745000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.375000 0.420000 0.985000 0.490000 ;
        RECT 0.375000 0.490000 0.510000 0.660000 ;
        RECT 0.915000 0.490000 0.985000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.07755 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2652 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185000 0.525000 0.255000 0.700000 ;
        RECT 0.185000 0.700000 0.320000 0.770000 ;
        RECT 0.185000 0.770000 1.200000 0.840000 ;
        RECT 1.130000 0.525000 1.200000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1099 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4095 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.415000 0.260000 1.485000 0.560000 ;
        RECT 1.415000 0.560000 1.860000 0.700000 ;
        RECT 1.415000 0.700000 1.485000 1.250000 ;
        RECT 1.790000 0.700000 1.860000 1.250000 ;
        RECT 1.790000 0.260000 1.860000 0.560000 ;
    END
    ANTENNADIFFAREA 0.297825 ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5941 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 1.210000 1.045000 1.280000 1.315000 ;
        RECT 0.075000 1.035000 0.145000 1.315000 ;
        RECT 1.595000 1.035000 1.665000 1.315000 ;
        RECT 1.975000 1.035000 2.045000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.075000 0.085000 0.145000 0.335000 ;
        RECT 0.450000 0.085000 0.520000 0.195000 ;
        RECT 0.830000 0.085000 0.900000 0.195000 ;
        RECT 1.210000 0.085000 1.280000 0.195000 ;
        RECT 1.595000 0.085000 1.665000 0.335000 ;
        RECT 1.975000 0.085000 2.045000 0.335000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.650000 0.980000 0.720000 1.250000 ;
      RECT 0.650000 0.910000 1.350000 0.980000 ;
      RECT 1.280000 0.330000 1.350000 0.910000 ;
      RECT 0.235000 0.260000 1.350000 0.330000 ;
  END
END OR3_X4

MACRO OR4_X1
  CLASS CORE ;
  FOREIGN OR4_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.760000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.990000 0.150000 1.080000 1.240000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0981 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3068 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.795000 0.965000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.285000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.900000 0.115000 1.240000 ;
      RECT 0.045000 0.830000 0.920000 0.900000 ;
      RECT 0.850000 0.420000 0.920000 0.830000 ;
      RECT 0.235000 0.350000 0.920000 0.420000 ;
      RECT 0.235000 0.150000 0.305000 0.350000 ;
      RECT 0.605000 0.150000 0.675000 0.350000 ;
  END
END OR4_X1

MACRO OR4_X2
  CLASS CORE ;
  FOREIGN OR4_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.760000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.150000 1.080000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
        RECT 1.175000 0.975000 1.245000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.285000 ;
        RECT 1.175000 0.085000 1.245000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.910000 0.115000 1.250000 ;
      RECT 0.045000 0.840000 0.925000 0.910000 ;
      RECT 0.855000 0.425000 0.925000 0.840000 ;
      RECT 0.235000 0.355000 0.925000 0.425000 ;
      RECT 0.235000 0.150000 0.305000 0.355000 ;
      RECT 0.605000 0.150000 0.675000 0.355000 ;
  END
END OR4_X2

MACRO OR4_X4
  CLASS CORE ;
  FOREIGN OR4_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.505000 0.390000 1.140000 0.460000 ;
        RECT 0.505000 0.460000 0.575000 0.660000 ;
        RECT 1.010000 0.460000 1.140000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08445 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2873 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
        RECT 0.310000 0.700000 0.380000 0.770000 ;
        RECT 0.310000 0.770000 1.330000 0.840000 ;
        RECT 1.260000 0.525000 1.330000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1162 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4264 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
        RECT 0.115000 0.700000 0.185000 0.905000 ;
        RECT 0.115000 0.905000 1.520000 0.975000 ;
        RECT 1.450000 0.525000 1.520000 0.905000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.161175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5954 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.755000 0.150000 1.825000 0.560000 ;
        RECT 1.755000 0.560000 2.200000 0.700000 ;
        RECT 1.755000 0.700000 1.825000 1.250000 ;
        RECT 2.130000 0.700000 2.200000 1.250000 ;
        RECT 2.130000 0.150000 2.200000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6513 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 1.555000 1.205000 1.625000 1.315000 ;
        RECT 0.040000 1.045000 0.110000 1.315000 ;
        RECT 1.935000 1.045000 2.005000 1.315000 ;
        RECT 2.315000 1.045000 2.385000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.400000 ;
        RECT 0.385000 0.085000 0.520000 0.160000 ;
        RECT 0.765000 0.085000 0.900000 0.160000 ;
        RECT 1.145000 0.085000 1.280000 0.160000 ;
        RECT 1.525000 0.085000 1.660000 0.325000 ;
        RECT 1.905000 0.085000 2.040000 0.365000 ;
        RECT 2.315000 0.085000 2.385000 0.400000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.770000 1.040000 1.685000 1.110000 ;
      RECT 1.615000 0.460000 1.685000 1.040000 ;
      RECT 1.370000 0.390000 1.685000 0.460000 ;
      RECT 1.370000 0.295000 1.440000 0.390000 ;
      RECT 0.235000 0.225000 1.440000 0.295000 ;
      RECT 0.235000 0.295000 0.305000 0.425000 ;
      RECT 0.235000 0.150000 0.305000 0.225000 ;
      RECT 1.370000 0.150000 1.440000 0.225000 ;
  END
END OR4_X4

MACRO SDFFRS_X1
  CLASS CORE ;
  FOREIGN SDFFRS_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 5.51 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.070000 0.765000 5.260000 0.980000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.04085 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1053 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.525000 0.920000 0.700000 ;
    END
    ANTENNAGATEAREA 0.0615 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.0615 LAYER metal2 ;
    ANTENNAGATEAREA 0.0615 LAYER metal3 ;
    ANTENNAGATEAREA 0.0615 LAYER metal4 ;
    ANTENNAGATEAREA 0.0615 LAYER metal5 ;
    ANTENNAGATEAREA 0.0615 LAYER metal6 ;
    ANTENNAGATEAREA 0.0615 LAYER metal7 ;
    ANTENNAGATEAREA 0.0615 LAYER metal8 ;
    ANTENNAGATEAREA 0.0615 LAYER metal9 ;
    ANTENNAGATEAREA 0.0615 LAYER metal10 ;
  END RN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.760000 0.390000 5.335000 0.460000 ;
        RECT 4.760000 0.460000 4.830000 0.765000 ;
        RECT 5.190000 0.460000 5.335000 0.560000 ;
        RECT 4.760000 0.765000 5.005000 0.835000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3367 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.560000 0.695000 4.690000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01885 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.110000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.575000 0.700000 1.670000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0133 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0611 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.045000 0.260000 0.130000 1.105000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.071825 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2418 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.360000 0.510000 0.800000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0374 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1365 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 5.510000 1.485000 ;
        RECT 0.195000 1.180000 0.330000 1.315000 ;
        RECT 4.415000 1.130000 4.550000 1.315000 ;
        RECT 0.925000 1.105000 1.060000 1.315000 ;
        RECT 1.305000 1.105000 1.440000 1.315000 ;
        RECT 5.175000 1.095000 5.310000 1.315000 ;
        RECT 0.545000 1.035000 0.680000 1.315000 ;
        RECT 3.585000 1.030000 3.720000 1.315000 ;
        RECT 2.665000 0.990000 2.800000 1.315000 ;
        RECT 3.045000 0.865000 3.180000 1.315000 ;
        RECT 1.945000 0.830000 2.015000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 5.510000 0.085000 ;
        RECT 0.195000 0.085000 0.330000 0.160000 ;
        RECT 0.920000 0.085000 1.055000 0.285000 ;
        RECT 1.755000 0.085000 1.825000 0.320000 ;
        RECT 2.665000 0.085000 2.800000 0.285000 ;
        RECT 3.400000 0.085000 3.535000 0.285000 ;
        RECT 4.415000 0.085000 4.550000 0.225000 ;
        RECT 5.175000 0.085000 5.310000 0.225000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.195000 0.900000 0.865000 0.970000 ;
      RECT 0.195000 0.295000 0.265000 0.900000 ;
      RECT 0.195000 0.225000 0.680000 0.295000 ;
      RECT 1.585000 1.165000 1.815000 1.235000 ;
      RECT 1.585000 0.975000 1.655000 1.165000 ;
      RECT 1.280000 0.905000 1.655000 0.975000 ;
      RECT 1.280000 0.480000 1.350000 0.905000 ;
      RECT 1.280000 0.410000 1.555000 0.480000 ;
      RECT 1.485000 0.285000 1.555000 0.410000 ;
      RECT 1.145000 0.835000 1.215000 1.105000 ;
      RECT 0.610000 0.765000 1.215000 0.835000 ;
      RECT 0.610000 0.460000 0.680000 0.765000 ;
      RECT 0.610000 0.390000 1.190000 0.460000 ;
      RECT 1.120000 0.320000 1.190000 0.390000 ;
      RECT 1.120000 0.250000 1.400000 0.320000 ;
      RECT 1.330000 0.220000 1.400000 0.250000 ;
      RECT 1.330000 0.150000 1.690000 0.220000 ;
      RECT 1.620000 0.220000 1.690000 0.385000 ;
      RECT 1.620000 0.385000 2.150000 0.455000 ;
      RECT 1.755000 0.765000 1.825000 0.965000 ;
      RECT 1.755000 0.695000 2.195000 0.765000 ;
      RECT 2.125000 0.765000 2.195000 0.965000 ;
      RECT 2.315000 0.625000 2.385000 0.965000 ;
      RECT 1.415000 0.555000 2.385000 0.625000 ;
      RECT 2.315000 0.200000 2.385000 0.555000 ;
      RECT 2.615000 0.755000 2.990000 0.825000 ;
      RECT 2.615000 0.555000 2.685000 0.755000 ;
      RECT 2.615000 0.485000 3.800000 0.555000 ;
      RECT 3.045000 0.295000 3.180000 0.485000 ;
      RECT 3.435000 0.965000 3.505000 1.115000 ;
      RECT 3.435000 0.895000 3.875000 0.965000 ;
      RECT 3.805000 0.965000 3.875000 1.115000 ;
      RECT 4.075000 0.690000 4.145000 1.115000 ;
      RECT 2.750000 0.620000 4.145000 0.690000 ;
      RECT 4.000000 0.295000 4.145000 0.620000 ;
      RECT 3.940000 1.180000 4.280000 1.250000 ;
      RECT 3.940000 0.830000 4.010000 1.180000 ;
      RECT 4.210000 0.230000 4.280000 1.180000 ;
      RECT 3.270000 0.760000 4.010000 0.830000 ;
      RECT 3.865000 0.160000 4.280000 0.230000 ;
      RECT 3.270000 0.830000 3.340000 1.090000 ;
      RECT 3.865000 0.230000 3.935000 0.350000 ;
      RECT 3.265000 0.350000 3.935000 0.420000 ;
      RECT 3.865000 0.420000 3.935000 0.510000 ;
      RECT 3.265000 0.230000 3.335000 0.350000 ;
      RECT 2.910000 0.160000 3.335000 0.230000 ;
      RECT 2.910000 0.230000 2.980000 0.350000 ;
      RECT 2.455000 0.350000 2.980000 0.420000 ;
      RECT 2.455000 0.420000 2.525000 1.035000 ;
      RECT 2.180000 1.035000 2.525000 1.105000 ;
      RECT 4.370000 0.945000 4.930000 1.015000 ;
      RECT 4.370000 0.480000 4.440000 0.945000 ;
      RECT 4.370000 0.410000 4.685000 0.480000 ;
      RECT 4.615000 0.290000 4.685000 0.410000 ;
      RECT 4.615000 0.220000 4.930000 0.290000 ;
      RECT 5.400000 0.695000 5.470000 1.235000 ;
      RECT 4.900000 0.625000 5.470000 0.695000 ;
      RECT 4.900000 0.560000 4.975000 0.625000 ;
      RECT 5.400000 0.215000 5.470000 0.625000 ;
  END
END SDFFRS_X1

MACRO SDFFRS_X2
  CLASS CORE ;
  FOREIGN SDFFRS_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 5.89 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.495000 0.420000 5.640000 0.560000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.545000 1.165000 0.700000 ;
    END
    ANTENNAGATEAREA 0.075 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.024025 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.075 LAYER metal2 ;
    ANTENNAGATEAREA 0.075 LAYER metal3 ;
    ANTENNAGATEAREA 0.075 LAYER metal4 ;
    ANTENNAGATEAREA 0.075 LAYER metal5 ;
    ANTENNAGATEAREA 0.075 LAYER metal6 ;
    ANTENNAGATEAREA 0.075 LAYER metal7 ;
    ANTENNAGATEAREA 0.075 LAYER metal8 ;
    ANTENNAGATEAREA 0.075 LAYER metal9 ;
    ANTENNAGATEAREA 0.075 LAYER metal10 ;
  END RN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.135000 0.385000 5.205000 0.720000 ;
        RECT 5.135000 0.720000 5.700000 0.790000 ;
        RECT 5.570000 0.790000 5.700000 0.840000 ;
        RECT 5.570000 0.675000 5.700000 0.720000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.07535 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2769 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.925000 0.560000 5.070000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.365000 0.545000 1.460000 0.700000 ;
    END
    ANTENNAGATEAREA 0.04875 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.065 LAYER metal1 ;
    ANTENNAGATEAREA 0.04875 LAYER metal2 ;
    ANTENNAGATEAREA 0.04875 LAYER metal3 ;
    ANTENNAGATEAREA 0.04875 LAYER metal4 ;
    ANTENNAGATEAREA 0.04875 LAYER metal5 ;
    ANTENNAGATEAREA 0.04875 LAYER metal6 ;
    ANTENNAGATEAREA 0.04875 LAYER metal7 ;
    ANTENNAGATEAREA 0.04875 LAYER metal8 ;
    ANTENNAGATEAREA 0.04875 LAYER metal9 ;
    ANTENNAGATEAREA 0.04875 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.900000 0.175000 2.065000 0.245000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0611 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.240000 0.150000 0.320000 1.125000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.078 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2743 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.600000 0.435000 0.735000 0.900000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.062775 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.156 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 5.890000 1.485000 ;
        RECT 5.540000 1.195000 5.675000 1.315000 ;
        RECT 1.180000 1.120000 1.315000 1.315000 ;
        RECT 1.640000 1.115000 1.775000 1.315000 ;
        RECT 0.410000 1.100000 0.545000 1.315000 ;
        RECT 0.790000 1.100000 0.925000 1.315000 ;
        RECT 3.950000 1.090000 4.085000 1.315000 ;
        RECT 4.780000 1.090000 4.915000 1.315000 ;
        RECT 3.040000 0.985000 3.175000 1.315000 ;
        RECT 3.420000 0.985000 3.555000 1.315000 ;
        RECT 2.285000 0.965000 2.420000 1.315000 ;
        RECT 0.065000 0.850000 0.135000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 5.890000 0.085000 ;
        RECT 0.065000 0.085000 0.135000 0.410000 ;
        RECT 0.410000 0.085000 0.545000 0.160000 ;
        RECT 0.790000 0.085000 0.925000 0.160000 ;
        RECT 1.700000 0.085000 1.835000 0.285000 ;
        RECT 2.130000 0.085000 2.200000 0.320000 ;
        RECT 3.040000 0.085000 3.175000 0.285000 ;
        RECT 3.760000 0.085000 3.895000 0.285000 ;
        RECT 4.810000 0.085000 4.880000 0.270000 ;
        RECT 5.540000 0.085000 5.675000 0.180000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.390000 0.965000 1.120000 1.035000 ;
      RECT 0.390000 0.300000 0.460000 0.965000 ;
      RECT 0.390000 0.230000 1.305000 0.300000 ;
      RECT 1.840000 1.160000 2.220000 1.230000 ;
      RECT 1.840000 1.045000 1.910000 1.160000 ;
      RECT 1.395000 0.975000 1.910000 1.045000 ;
      RECT 1.395000 0.835000 1.465000 0.975000 ;
      RECT 0.870000 0.765000 1.465000 0.835000 ;
      RECT 0.870000 0.480000 0.940000 0.765000 ;
      RECT 0.870000 0.410000 1.460000 0.480000 ;
      RECT 2.130000 0.900000 2.200000 1.050000 ;
      RECT 2.130000 0.830000 2.570000 0.900000 ;
      RECT 2.500000 0.900000 2.570000 1.050000 ;
      RECT 1.530000 0.840000 2.040000 0.910000 ;
      RECT 1.970000 0.755000 2.040000 0.840000 ;
      RECT 1.530000 0.420000 1.600000 0.840000 ;
      RECT 1.970000 0.685000 2.635000 0.755000 ;
      RECT 1.530000 0.350000 2.040000 0.420000 ;
      RECT 2.565000 0.620000 2.635000 0.685000 ;
      RECT 1.665000 0.555000 1.735000 0.680000 ;
      RECT 1.665000 0.485000 2.770000 0.555000 ;
      RECT 2.700000 0.555000 2.770000 1.050000 ;
      RECT 2.700000 0.200000 2.770000 0.485000 ;
      RECT 2.990000 0.765000 3.370000 0.835000 ;
      RECT 2.990000 0.560000 3.060000 0.765000 ;
      RECT 2.990000 0.490000 4.170000 0.560000 ;
      RECT 2.990000 0.485000 3.525000 0.490000 ;
      RECT 3.455000 0.320000 3.525000 0.485000 ;
      RECT 3.800000 1.025000 3.870000 1.175000 ;
      RECT 3.800000 0.955000 4.240000 1.025000 ;
      RECT 4.170000 1.025000 4.240000 1.175000 ;
      RECT 4.440000 0.695000 4.510000 1.090000 ;
      RECT 3.125000 0.625000 4.510000 0.695000 ;
      RECT 4.405000 0.355000 4.475000 0.625000 ;
      RECT 4.405000 0.285000 4.540000 0.355000 ;
      RECT 2.555000 1.115000 2.915000 1.185000 ;
      RECT 2.845000 0.420000 2.915000 1.115000 ;
      RECT 2.845000 0.350000 3.390000 0.420000 ;
      RECT 3.320000 0.220000 3.390000 0.350000 ;
      RECT 3.320000 0.150000 3.680000 0.220000 ;
      RECT 3.610000 0.220000 3.680000 0.355000 ;
      RECT 3.610000 0.355000 4.340000 0.425000 ;
      RECT 4.270000 0.220000 4.340000 0.355000 ;
      RECT 4.270000 0.150000 4.675000 0.220000 ;
      RECT 4.605000 0.220000 4.675000 0.690000 ;
      RECT 4.575000 0.690000 4.675000 0.825000 ;
      RECT 4.605000 0.825000 4.675000 1.155000 ;
      RECT 4.305000 1.155000 4.675000 1.225000 ;
      RECT 4.305000 0.835000 4.375000 1.155000 ;
      RECT 3.615000 0.765000 4.375000 0.835000 ;
      RECT 4.740000 0.950000 5.295000 1.020000 ;
      RECT 4.740000 0.445000 4.810000 0.950000 ;
      RECT 4.740000 0.375000 5.045000 0.445000 ;
      RECT 4.975000 0.235000 5.045000 0.375000 ;
      RECT 4.975000 0.165000 5.295000 0.235000 ;
      RECT 5.270000 0.565000 5.410000 0.635000 ;
      RECT 5.340000 0.355000 5.410000 0.565000 ;
      RECT 5.340000 0.285000 5.835000 0.355000 ;
      RECT 5.765000 0.355000 5.835000 1.090000 ;
      RECT 5.765000 0.150000 5.835000 0.285000 ;
  END
END SDFFRS_X2

MACRO SDFFR_X1
  CLASS CORE ;
  FOREIGN SDFFR_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.75 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.240000 0.560000 4.365000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.840000 0.925000 0.980000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0147 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END RN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.105000 0.565000 4.175000 0.770000 ;
        RECT 4.105000 0.770000 4.530000 0.840000 ;
        RECT 4.430000 0.560000 4.530000 0.770000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0651 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2366 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.670000 0.655000 3.765000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.017575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.770000 0.660000 1.995000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0405 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1053 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.435000 0.185000 0.510000 1.015000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.06225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2353 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.185000 0.130000 1.065000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0616 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.247 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.750000 1.485000 ;
        RECT 0.210000 1.240000 0.345000 1.315000 ;
        RECT 0.740000 1.240000 0.875000 1.315000 ;
        RECT 1.150000 1.205000 1.220000 1.315000 ;
        RECT 3.270000 1.080000 3.340000 1.315000 ;
        RECT 3.640000 1.080000 3.710000 1.315000 ;
        RECT 1.840000 1.060000 1.975000 1.315000 ;
        RECT 4.400000 1.045000 4.470000 1.315000 ;
        RECT 2.400000 0.995000 2.470000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.750000 0.085000 ;
        RECT 0.240000 0.085000 0.310000 0.460000 ;
        RECT 0.770000 0.085000 0.840000 0.320000 ;
        RECT 1.710000 0.085000 1.845000 0.285000 ;
        RECT 2.270000 0.085000 2.340000 0.425000 ;
        RECT 3.110000 0.085000 3.180000 0.320000 ;
        RECT 3.640000 0.085000 3.710000 0.320000 ;
        RECT 4.400000 0.085000 4.470000 0.320000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.585000 1.150000 0.655000 1.240000 ;
      RECT 0.195000 1.080000 0.655000 1.150000 ;
      RECT 0.195000 0.525000 0.265000 1.080000 ;
      RECT 0.585000 0.460000 0.655000 1.080000 ;
      RECT 0.585000 0.390000 1.075000 0.460000 ;
      RECT 1.005000 0.460000 1.075000 0.635000 ;
      RECT 0.585000 0.185000 0.655000 0.390000 ;
      RECT 0.935000 1.045000 1.410000 1.115000 ;
      RECT 1.490000 0.975000 1.560000 1.040000 ;
      RECT 1.140000 0.905000 1.560000 0.975000 ;
      RECT 1.140000 0.775000 1.210000 0.905000 ;
      RECT 0.720000 0.705000 1.210000 0.775000 ;
      RECT 0.720000 0.525000 0.790000 0.705000 ;
      RECT 1.140000 0.285000 1.210000 0.705000 ;
      RECT 1.140000 0.215000 1.460000 0.285000 ;
      RECT 1.545000 1.180000 1.695000 1.250000 ;
      RECT 1.625000 0.975000 1.695000 1.180000 ;
      RECT 1.625000 0.905000 2.135000 0.975000 ;
      RECT 2.065000 0.975000 2.135000 1.065000 ;
      RECT 1.625000 0.835000 1.695000 0.905000 ;
      RECT 2.065000 0.790000 2.135000 0.905000 ;
      RECT 1.280000 0.765000 1.695000 0.835000 ;
      RECT 2.065000 0.655000 2.260000 0.790000 ;
      RECT 1.280000 0.420000 1.350000 0.765000 ;
      RECT 1.280000 0.350000 2.000000 0.420000 ;
      RECT 1.930000 0.185000 2.000000 0.350000 ;
      RECT 2.220000 0.925000 2.290000 1.130000 ;
      RECT 2.220000 0.855000 2.405000 0.925000 ;
      RECT 2.335000 0.560000 2.405000 0.855000 ;
      RECT 1.430000 0.490000 2.475000 0.560000 ;
      RECT 1.430000 0.560000 1.500000 0.700000 ;
      RECT 2.405000 0.240000 2.475000 0.490000 ;
      RECT 2.090000 0.185000 2.160000 0.490000 ;
      RECT 2.405000 0.170000 2.920000 0.240000 ;
      RECT 2.850000 0.240000 2.920000 0.835000 ;
      RECT 2.690000 1.015000 3.065000 1.085000 ;
      RECT 2.995000 0.880000 3.065000 1.015000 ;
      RECT 2.690000 0.305000 2.760000 1.015000 ;
      RECT 2.995000 0.810000 3.450000 0.880000 ;
      RECT 2.540000 1.180000 3.205000 1.250000 ;
      RECT 3.135000 1.015000 3.205000 1.180000 ;
      RECT 2.540000 0.505000 2.610000 1.180000 ;
      RECT 3.135000 0.945000 3.585000 1.015000 ;
      RECT 3.450000 1.015000 3.520000 1.200000 ;
      RECT 3.515000 0.725000 3.585000 0.945000 ;
      RECT 2.985000 0.655000 3.585000 0.725000 ;
      RECT 2.985000 0.455000 3.055000 0.655000 ;
      RECT 2.985000 0.385000 3.335000 0.455000 ;
      RECT 3.265000 0.185000 3.335000 0.385000 ;
      RECT 3.830000 1.040000 4.125000 1.110000 ;
      RECT 3.830000 0.590000 3.900000 1.040000 ;
      RECT 3.120000 0.520000 3.900000 0.590000 ;
      RECT 3.830000 0.290000 3.900000 0.520000 ;
      RECT 3.830000 0.220000 4.125000 0.290000 ;
      RECT 4.595000 0.975000 4.665000 1.220000 ;
      RECT 3.965000 0.905000 4.665000 0.975000 ;
      RECT 3.965000 0.715000 4.035000 0.905000 ;
      RECT 4.595000 0.485000 4.665000 0.905000 ;
      RECT 4.100000 0.415000 4.665000 0.485000 ;
      RECT 4.595000 0.185000 4.665000 0.415000 ;
  END
END SDFFR_X1

MACRO SDFFR_X2
  CLASS CORE ;
  FOREIGN SDFFR_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.565000 0.420000 4.690000 0.625000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.025625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145000 0.840000 1.270000 0.980000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END RN

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.345000 0.565000 4.415000 0.700000 ;
        RECT 4.345000 0.700000 4.765000 0.845000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.07035 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.182 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.860000 0.670000 4.005000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02465 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0819 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.145000 0.695000 2.280000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.019575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.395000 0.510000 1.005000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.05185 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1807 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.795000 0.395000 0.865000 0.560000 ;
        RECT 0.795000 0.560000 0.890000 1.005000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.053825 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1833 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.940000 1.485000 ;
        RECT 0.575000 1.240000 0.710000 1.315000 ;
        RECT 0.225000 1.205000 0.295000 1.315000 ;
        RECT 0.985000 1.205000 1.055000 1.315000 ;
        RECT 1.370000 1.205000 1.440000 1.315000 ;
        RECT 3.460000 1.115000 3.595000 1.315000 ;
        RECT 3.875000 1.080000 3.945000 1.315000 ;
        RECT 2.060000 1.060000 2.195000 1.315000 ;
        RECT 4.635000 1.045000 4.705000 1.315000 ;
        RECT 2.660000 0.995000 2.730000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.940000 0.085000 ;
        RECT 0.195000 0.085000 0.330000 0.160000 ;
        RECT 0.575000 0.085000 0.710000 0.160000 ;
        RECT 1.065000 0.085000 1.135000 0.320000 ;
        RECT 2.005000 0.085000 2.075000 0.320000 ;
        RECT 2.535000 0.085000 2.605000 0.420000 ;
        RECT 3.295000 0.085000 3.365000 0.320000 ;
        RECT 3.875000 0.085000 3.945000 0.320000 ;
        RECT 4.635000 0.085000 4.705000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 1.070000 1.080000 1.140000 ;
      RECT 1.010000 0.775000 1.080000 1.070000 ;
      RECT 0.660000 0.525000 0.730000 1.070000 ;
      RECT 0.045000 0.260000 0.115000 1.070000 ;
      RECT 1.010000 0.640000 1.360000 0.775000 ;
      RECT 1.155000 1.115000 1.290000 1.250000 ;
      RECT 1.155000 1.045000 1.630000 1.115000 ;
      RECT 1.425000 0.885000 1.815000 0.955000 ;
      RECT 1.425000 0.455000 1.495000 0.885000 ;
      RECT 0.930000 0.385000 1.495000 0.455000 ;
      RECT 1.425000 0.335000 1.495000 0.385000 ;
      RECT 0.930000 0.330000 1.000000 0.385000 ;
      RECT 1.425000 0.265000 1.730000 0.335000 ;
      RECT 0.290000 0.260000 1.000000 0.330000 ;
      RECT 0.290000 0.330000 0.360000 0.660000 ;
      RECT 1.790000 1.180000 1.950000 1.250000 ;
      RECT 1.880000 0.985000 1.950000 1.180000 ;
      RECT 1.880000 0.915000 2.415000 0.985000 ;
      RECT 1.880000 0.820000 1.950000 0.915000 ;
      RECT 2.345000 0.750000 2.415000 0.915000 ;
      RECT 1.560000 0.750000 1.950000 0.820000 ;
      RECT 2.345000 0.680000 2.560000 0.750000 ;
      RECT 1.560000 0.480000 1.630000 0.750000 ;
      RECT 1.560000 0.410000 2.265000 0.480000 ;
      RECT 2.195000 0.260000 2.265000 0.410000 ;
      RECT 2.480000 0.885000 2.550000 1.090000 ;
      RECT 2.480000 0.815000 2.740000 0.885000 ;
      RECT 2.670000 0.615000 2.740000 0.815000 ;
      RECT 1.715000 0.545000 2.740000 0.615000 ;
      RECT 1.715000 0.615000 1.785000 0.685000 ;
      RECT 2.350000 0.285000 2.420000 0.545000 ;
      RECT 2.670000 0.235000 2.740000 0.545000 ;
      RECT 2.670000 0.165000 3.220000 0.235000 ;
      RECT 3.150000 0.235000 3.220000 0.775000 ;
      RECT 3.040000 0.915000 3.110000 1.115000 ;
      RECT 2.955000 0.910000 3.110000 0.915000 ;
      RECT 2.955000 0.840000 3.625000 0.910000 ;
      RECT 2.955000 0.400000 3.025000 0.840000 ;
      RECT 2.890000 0.330000 3.025000 0.400000 ;
      RECT 2.805000 1.180000 3.255000 1.250000 ;
      RECT 3.185000 1.045000 3.255000 1.180000 ;
      RECT 2.805000 0.500000 2.875000 1.180000 ;
      RECT 3.185000 0.975000 3.760000 1.045000 ;
      RECT 3.690000 1.045000 3.760000 1.200000 ;
      RECT 3.690000 0.725000 3.760000 0.975000 ;
      RECT 3.285000 0.655000 3.760000 0.725000 ;
      RECT 3.285000 0.455000 3.355000 0.655000 ;
      RECT 3.285000 0.385000 3.570000 0.455000 ;
      RECT 3.500000 0.200000 3.570000 0.385000 ;
      RECT 4.070000 1.045000 4.360000 1.115000 ;
      RECT 4.070000 0.590000 4.140000 1.045000 ;
      RECT 3.420000 0.520000 4.140000 0.590000 ;
      RECT 4.070000 0.300000 4.140000 0.520000 ;
      RECT 4.070000 0.230000 4.360000 0.300000 ;
      RECT 4.830000 0.980000 4.900000 1.220000 ;
      RECT 4.205000 0.910000 4.900000 0.980000 ;
      RECT 4.205000 0.715000 4.275000 0.910000 ;
      RECT 4.830000 0.355000 4.900000 0.910000 ;
      RECT 4.425000 0.285000 4.900000 0.355000 ;
      RECT 4.425000 0.355000 4.495000 0.415000 ;
      RECT 4.830000 0.195000 4.900000 0.285000 ;
      RECT 4.360000 0.415000 4.495000 0.485000 ;
  END
END SDFFR_X2

MACRO SDFFS_X1
  CLASS CORE ;
  FOREIGN SDFFS_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.75 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.550000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0195 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.550000 0.185000 0.765000 ;
        RECT 0.060000 0.765000 0.570000 0.835000 ;
        RECT 0.500000 0.550000 0.570000 0.765000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.077625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2626 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.910000 0.420000 1.080000 0.560000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.840000 0.420000 3.930000 0.575000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01395 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.785000 1.115000 0.980000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.020475 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.240000 0.980000 4.335000 1.250000 ;
        RECT 4.265000 0.400000 4.335000 0.980000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.06625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2457 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.620000 0.980000 4.705000 1.250000 ;
        RECT 4.635000 0.150000 4.705000 0.980000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.08105 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.750000 1.485000 ;
        RECT 2.300000 1.155000 2.370000 1.315000 ;
        RECT 2.830000 1.070000 2.900000 1.315000 ;
        RECT 3.735000 1.070000 3.805000 1.315000 ;
        RECT 0.985000 1.045000 1.055000 1.315000 ;
        RECT 1.520000 1.040000 1.590000 1.315000 ;
        RECT 0.225000 1.035000 0.295000 1.315000 ;
        RECT 4.105000 0.975000 4.175000 1.315000 ;
        RECT 4.445000 0.975000 4.515000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.750000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.985000 0.085000 1.055000 0.285000 ;
        RECT 1.490000 0.085000 1.625000 0.215000 ;
        RECT 2.485000 0.085000 2.555000 0.370000 ;
        RECT 2.805000 0.085000 2.940000 0.285000 ;
        RECT 3.735000 0.085000 3.805000 0.320000 ;
        RECT 4.445000 0.085000 4.515000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.970000 0.115000 1.250000 ;
      RECT 0.045000 0.900000 0.765000 0.970000 ;
      RECT 0.635000 0.835000 0.765000 0.900000 ;
      RECT 0.635000 0.485000 0.705000 0.835000 ;
      RECT 0.045000 0.415000 0.705000 0.485000 ;
      RECT 0.045000 0.150000 0.115000 0.415000 ;
      RECT 0.580000 1.105000 0.715000 1.240000 ;
      RECT 0.580000 1.035000 0.900000 1.105000 ;
      RECT 0.830000 0.695000 0.900000 1.035000 ;
      RECT 0.775000 0.625000 1.540000 0.695000 ;
      RECT 0.775000 0.285000 0.845000 0.625000 ;
      RECT 0.615000 0.150000 0.845000 0.285000 ;
      RECT 1.180000 0.840000 1.250000 1.250000 ;
      RECT 1.180000 0.770000 1.675000 0.840000 ;
      RECT 1.605000 0.670000 1.675000 0.770000 ;
      RECT 1.605000 0.600000 1.890000 0.670000 ;
      RECT 1.605000 0.485000 1.675000 0.600000 ;
      RECT 1.180000 0.415000 1.675000 0.485000 ;
      RECT 1.180000 0.150000 1.250000 0.415000 ;
      RECT 2.070000 1.170000 2.205000 1.240000 ;
      RECT 2.135000 1.090000 2.205000 1.170000 ;
      RECT 2.135000 1.020000 2.525000 1.090000 ;
      RECT 2.455000 1.090000 2.525000 1.170000 ;
      RECT 2.455000 1.170000 2.590000 1.240000 ;
      RECT 1.870000 1.170000 2.005000 1.240000 ;
      RECT 1.935000 0.950000 2.005000 1.170000 ;
      RECT 1.935000 0.880000 2.160000 0.950000 ;
      RECT 2.090000 0.735000 2.160000 0.880000 ;
      RECT 2.090000 0.665000 2.945000 0.735000 ;
      RECT 2.090000 0.355000 2.160000 0.665000 ;
      RECT 1.875000 0.285000 2.160000 0.355000 ;
      RECT 1.340000 0.975000 1.410000 1.250000 ;
      RECT 1.340000 0.905000 1.865000 0.975000 ;
      RECT 1.795000 0.810000 1.865000 0.905000 ;
      RECT 1.795000 0.740000 2.025000 0.810000 ;
      RECT 1.955000 0.490000 2.025000 0.740000 ;
      RECT 1.740000 0.420000 2.025000 0.490000 ;
      RECT 1.740000 0.350000 1.810000 0.420000 ;
      RECT 1.340000 0.280000 1.810000 0.350000 ;
      RECT 1.740000 0.220000 1.810000 0.280000 ;
      RECT 1.340000 0.150000 1.410000 0.280000 ;
      RECT 1.740000 0.150000 2.295000 0.220000 ;
      RECT 2.225000 0.220000 2.295000 0.485000 ;
      RECT 2.225000 0.485000 3.355000 0.555000 ;
      RECT 3.285000 0.555000 3.355000 0.860000 ;
      RECT 2.615000 0.930000 3.490000 1.000000 ;
      RECT 2.615000 0.875000 2.685000 0.930000 ;
      RECT 3.420000 0.420000 3.490000 0.930000 ;
      RECT 2.225000 0.805000 2.685000 0.875000 ;
      RECT 2.650000 0.350000 3.490000 0.420000 ;
      RECT 2.650000 0.200000 2.720000 0.350000 ;
      RECT 3.255000 1.100000 3.625000 1.170000 ;
      RECT 3.555000 0.710000 3.625000 1.100000 ;
      RECT 3.555000 0.640000 4.065000 0.710000 ;
      RECT 3.995000 0.525000 4.065000 0.640000 ;
      RECT 3.555000 0.285000 3.625000 0.640000 ;
      RECT 3.250000 0.215000 3.625000 0.285000 ;
      RECT 3.915000 0.915000 3.985000 1.250000 ;
      RECT 3.690000 0.845000 3.985000 0.915000 ;
      RECT 3.690000 0.775000 4.200000 0.845000 ;
      RECT 4.130000 0.335000 4.200000 0.775000 ;
      RECT 4.075000 0.265000 4.565000 0.335000 ;
      RECT 4.495000 0.335000 4.565000 0.660000 ;
  END
END SDFFS_X1

MACRO SDFFS_X2
  CLASS CORE ;
  FOREIGN SDFFS_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 5.13 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.670000 0.375000 0.840000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.795000 0.185000 0.910000 ;
        RECT 0.060000 0.910000 0.595000 0.980000 ;
        RECT 0.525000 0.670000 0.595000 0.910000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.068625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.965000 0.420000 1.080000 0.640000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0253 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0871 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.420000 0.425000 2.980000 0.495000 ;
        RECT 2.910000 0.350000 2.980000 0.425000 ;
        RECT 2.910000 0.280000 3.410000 0.350000 ;
        RECT 3.340000 0.350000 3.410000 0.560000 ;
        RECT 3.340000 0.560000 4.030000 0.630000 ;
    END
    ANTENNAGATEAREA 0.06125 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.14245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5473 LAYER metal1 ;
    ANTENNAGATEAREA 0.06125 LAYER metal2 ;
    ANTENNAGATEAREA 0.06125 LAYER metal3 ;
    ANTENNAGATEAREA 0.06125 LAYER metal4 ;
    ANTENNAGATEAREA 0.06125 LAYER metal5 ;
    ANTENNAGATEAREA 0.06125 LAYER metal6 ;
    ANTENNAGATEAREA 0.06125 LAYER metal7 ;
    ANTENNAGATEAREA 0.06125 LAYER metal8 ;
    ANTENNAGATEAREA 0.06125 LAYER metal9 ;
    ANTENNAGATEAREA 0.06125 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.840000 1.130000 0.980000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.430000 0.395000 4.500000 0.785000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0273 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1196 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.810000 0.395000 4.880000 0.785000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0273 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1196 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 5.130000 1.485000 ;
        RECT 0.195000 1.240000 0.330000 1.315000 ;
        RECT 1.505000 1.240000 1.640000 1.315000 ;
        RECT 2.265000 1.165000 2.400000 1.315000 ;
        RECT 3.825000 1.150000 3.960000 1.315000 ;
        RECT 4.200000 1.150000 4.335000 1.315000 ;
        RECT 4.580000 1.150000 4.715000 1.315000 ;
        RECT 4.990000 1.125000 5.060000 1.315000 ;
        RECT 3.510000 1.120000 3.580000 1.315000 ;
        RECT 0.990000 1.115000 1.060000 1.315000 ;
        RECT 2.640000 1.030000 2.710000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 5.130000 0.085000 ;
        RECT 0.200000 0.085000 0.335000 0.465000 ;
        RECT 0.960000 0.085000 1.095000 0.280000 ;
        RECT 1.510000 0.085000 1.645000 0.345000 ;
        RECT 2.475000 0.085000 2.610000 0.345000 ;
        RECT 3.475000 0.085000 3.610000 0.480000 ;
        RECT 4.200000 0.085000 4.335000 0.180000 ;
        RECT 4.580000 0.085000 4.715000 0.180000 ;
        RECT 4.990000 0.085000 5.060000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 1.115000 0.115000 1.250000 ;
      RECT 0.045000 1.045000 0.765000 1.115000 ;
      RECT 0.695000 0.605000 0.765000 1.045000 ;
      RECT 0.045000 0.535000 0.765000 0.605000 ;
      RECT 0.045000 0.380000 0.115000 0.535000 ;
      RECT 0.585000 1.180000 0.900000 1.250000 ;
      RECT 0.830000 0.775000 0.900000 1.180000 ;
      RECT 0.830000 0.705000 1.570000 0.775000 ;
      RECT 0.830000 0.420000 0.900000 0.705000 ;
      RECT 0.585000 0.350000 0.900000 0.420000 ;
      RECT 1.195000 0.940000 1.265000 1.250000 ;
      RECT 1.195000 0.870000 1.705000 0.940000 ;
      RECT 1.635000 0.695000 1.705000 0.870000 ;
      RECT 1.635000 0.630000 1.915000 0.695000 ;
      RECT 1.195000 0.625000 1.915000 0.630000 ;
      RECT 1.195000 0.560000 1.705000 0.625000 ;
      RECT 1.195000 0.315000 1.265000 0.560000 ;
      RECT 2.115000 1.100000 2.185000 1.250000 ;
      RECT 2.115000 1.030000 2.555000 1.100000 ;
      RECT 2.485000 1.100000 2.555000 1.250000 ;
      RECT 1.925000 0.965000 1.995000 1.250000 ;
      RECT 1.925000 0.895000 2.195000 0.965000 ;
      RECT 2.125000 0.765000 2.195000 0.895000 ;
      RECT 2.125000 0.695000 2.825000 0.765000 ;
      RECT 2.150000 0.360000 2.220000 0.695000 ;
      RECT 1.895000 0.290000 2.220000 0.360000 ;
      RECT 1.355000 1.175000 1.425000 1.250000 ;
      RECT 1.355000 1.105000 1.855000 1.175000 ;
      RECT 1.785000 0.830000 1.855000 1.105000 ;
      RECT 1.785000 0.760000 2.050000 0.830000 ;
      RECT 1.980000 0.575000 2.050000 0.760000 ;
      RECT 1.980000 0.495000 2.075000 0.575000 ;
      RECT 1.355000 0.425000 2.075000 0.495000 ;
      RECT 1.355000 0.360000 1.425000 0.425000 ;
      RECT 1.750000 0.225000 1.820000 0.425000 ;
      RECT 1.750000 0.155000 2.355000 0.225000 ;
      RECT 2.285000 0.225000 2.355000 0.560000 ;
      RECT 2.285000 0.560000 3.140000 0.630000 ;
      RECT 3.070000 0.630000 3.140000 0.845000 ;
      RECT 3.070000 0.845000 3.175000 0.980000 ;
      RECT 3.045000 1.045000 3.310000 1.115000 ;
      RECT 3.240000 0.765000 3.310000 1.045000 ;
      RECT 3.240000 0.760000 4.230000 0.765000 ;
      RECT 3.205000 0.695000 4.230000 0.760000 ;
      RECT 4.095000 0.560000 4.230000 0.695000 ;
      RECT 3.205000 0.485000 3.275000 0.695000 ;
      RECT 3.045000 0.415000 3.275000 0.485000 ;
      RECT 3.375000 0.850000 4.745000 0.920000 ;
      RECT 4.675000 0.525000 4.745000 0.850000 ;
      RECT 4.295000 0.485000 4.365000 0.850000 ;
      RECT 3.825000 0.415000 4.365000 0.485000 ;
      RECT 2.910000 1.180000 3.445000 1.250000 ;
      RECT 3.375000 1.055000 3.445000 1.180000 ;
      RECT 2.910000 0.965000 2.980000 1.180000 ;
      RECT 3.375000 0.985000 5.015000 1.055000 ;
      RECT 2.260000 0.830000 2.980000 0.965000 ;
      RECT 4.945000 0.330000 5.015000 0.985000 ;
      RECT 3.690000 0.260000 5.015000 0.330000 ;
      RECT 3.690000 0.330000 3.760000 0.495000 ;
  END
END SDFFS_X2

MACRO SDFF_X1
  CLASS CORE ;
  FOREIGN SDFF_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.37 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.975000 0.420000 4.125000 0.565000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.750000 0.590000 3.885000 0.700000 ;
        RECT 3.750000 0.700000 4.180000 0.770000 ;
        RECT 4.050000 0.770000 4.180000 0.840000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.05405 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1768 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.415000 0.525000 3.550000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.023625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.020000 0.420000 2.225000 0.580000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0328 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0949 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.150000 0.510000 0.785000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.04445 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1833 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.150000 0.135000 1.215000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.079875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2964 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.370000 1.485000 ;
        RECT 0.750000 1.165000 0.885000 1.315000 ;
        RECT 2.935000 1.080000 3.005000 1.315000 ;
        RECT 0.250000 1.040000 0.320000 1.315000 ;
        RECT 3.295000 1.040000 3.365000 1.315000 ;
        RECT 1.510000 0.975000 1.645000 1.315000 ;
        RECT 4.020000 0.975000 4.155000 1.315000 ;
        RECT 2.070000 0.940000 2.140000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.370000 0.085000 ;
        RECT 0.250000 0.085000 0.320000 0.425000 ;
        RECT 0.750000 0.085000 0.885000 0.285000 ;
        RECT 1.510000 0.085000 1.645000 0.285000 ;
        RECT 2.040000 0.085000 2.175000 0.285000 ;
        RECT 2.905000 0.085000 3.040000 0.190000 ;
        RECT 3.295000 0.085000 3.365000 0.195000 ;
        RECT 4.020000 0.085000 4.155000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.595000 0.955000 0.665000 1.215000 ;
      RECT 0.200000 0.885000 0.665000 0.955000 ;
      RECT 0.595000 0.865000 0.665000 0.885000 ;
      RECT 0.200000 0.510000 0.270000 0.885000 ;
      RECT 0.595000 0.730000 0.925000 0.865000 ;
      RECT 0.595000 0.150000 0.665000 0.730000 ;
      RECT 0.990000 1.150000 1.265000 1.220000 ;
      RECT 0.990000 0.660000 1.060000 1.150000 ;
      RECT 0.730000 0.525000 1.060000 0.660000 ;
      RECT 0.990000 0.300000 1.060000 0.525000 ;
      RECT 0.990000 0.230000 1.265000 0.300000 ;
      RECT 1.730000 0.910000 1.800000 1.215000 ;
      RECT 1.125000 0.840000 1.800000 0.910000 ;
      RECT 1.125000 0.545000 1.195000 0.840000 ;
      RECT 1.125000 0.475000 1.800000 0.545000 ;
      RECT 1.730000 0.320000 1.800000 0.475000 ;
      RECT 1.885000 0.750000 1.955000 1.090000 ;
      RECT 1.885000 0.720000 2.565000 0.750000 ;
      RECT 2.370000 0.750000 2.440000 0.950000 ;
      RECT 1.260000 0.680000 2.565000 0.720000 ;
      RECT 1.260000 0.650000 1.955000 0.680000 ;
      RECT 2.495000 0.350000 2.565000 0.680000 ;
      RECT 1.885000 0.200000 1.955000 0.650000 ;
      RECT 2.530000 0.975000 2.700000 1.045000 ;
      RECT 2.630000 0.460000 2.700000 0.975000 ;
      RECT 2.630000 0.325000 3.080000 0.460000 ;
      RECT 2.630000 0.285000 2.700000 0.325000 ;
      RECT 2.530000 0.215000 2.700000 0.285000 ;
      RECT 2.205000 1.140000 2.835000 1.210000 ;
      RECT 2.765000 0.990000 2.835000 1.140000 ;
      RECT 2.205000 0.815000 2.275000 1.140000 ;
      RECT 2.765000 0.920000 3.195000 0.990000 ;
      RECT 3.125000 0.990000 3.195000 1.215000 ;
      RECT 2.765000 0.615000 2.835000 0.920000 ;
      RECT 2.765000 0.545000 3.215000 0.615000 ;
      RECT 3.145000 0.150000 3.215000 0.545000 ;
      RECT 3.670000 0.975000 3.740000 1.215000 ;
      RECT 3.280000 0.905000 3.740000 0.975000 ;
      RECT 3.280000 0.830000 3.350000 0.905000 ;
      RECT 2.900000 0.695000 3.350000 0.830000 ;
      RECT 3.280000 0.355000 3.350000 0.695000 ;
      RECT 3.280000 0.285000 3.740000 0.355000 ;
      RECT 3.670000 0.150000 3.740000 0.285000 ;
      RECT 3.615000 0.520000 3.685000 0.840000 ;
      RECT 3.615000 0.450000 3.880000 0.520000 ;
      RECT 3.810000 0.350000 3.880000 0.450000 ;
      RECT 3.810000 0.280000 4.315000 0.350000 ;
      RECT 4.245000 0.350000 4.315000 1.215000 ;
      RECT 4.245000 0.150000 4.315000 0.280000 ;
  END
END SDFF_X1

MACRO SDFF_X2
  CLASS CORE ;
  FOREIGN SDFF_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.165000 0.420000 4.330000 0.560000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.950000 0.595000 4.020000 0.700000 ;
        RECT 3.950000 0.700000 4.355000 0.840000 ;
    END
    ANTENNAGATEAREA 0.05775 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.06405 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.169 LAYER metal1 ;
    ANTENNAGATEAREA 0.05775 LAYER metal2 ;
    ANTENNAGATEAREA 0.05775 LAYER metal3 ;
    ANTENNAGATEAREA 0.05775 LAYER metal4 ;
    ANTENNAGATEAREA 0.05775 LAYER metal5 ;
    ANTENNAGATEAREA 0.05775 LAYER metal6 ;
    ANTENNAGATEAREA 0.05775 LAYER metal7 ;
    ANTENNAGATEAREA 0.05775 LAYER metal8 ;
    ANTENNAGATEAREA 0.05775 LAYER metal9 ;
    ANTENNAGATEAREA 0.05775 LAYER metal10 ;
  END SE

  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.480000 0.420000 3.580000 0.560000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0624 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SI

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.225000 0.420000 2.410000 0.580000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0296 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0897 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.400000 0.510000 0.785000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.032725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1222 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805000 0.185000 0.890000 0.840000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.055675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1924 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.560000 1.485000 ;
        RECT 3.455000 1.240000 3.590000 1.315000 ;
        RECT 3.135000 1.080000 3.205000 1.315000 ;
        RECT 0.225000 1.040000 0.295000 1.315000 ;
        RECT 0.605000 1.040000 0.675000 1.315000 ;
        RECT 0.985000 1.040000 1.055000 1.315000 ;
        RECT 4.240000 0.965000 4.310000 1.315000 ;
        RECT 1.745000 0.940000 1.815000 1.315000 ;
        RECT 2.275000 0.910000 2.345000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.560000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.195000 ;
        RECT 0.605000 0.085000 0.675000 0.195000 ;
        RECT 0.985000 0.085000 1.055000 0.320000 ;
        RECT 1.745000 0.085000 1.815000 0.320000 ;
        RECT 2.275000 0.085000 2.345000 0.320000 ;
        RECT 3.065000 0.085000 3.200000 0.165000 ;
        RECT 3.485000 0.085000 3.555000 0.255000 ;
        RECT 4.210000 0.085000 4.345000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.335000 0.115000 1.185000 ;
      RECT 0.045000 0.265000 0.740000 0.335000 ;
      RECT 0.670000 0.335000 0.740000 0.660000 ;
      RECT 0.045000 0.185000 0.115000 0.265000 ;
      RECT 1.130000 1.055000 1.470000 1.125000 ;
      RECT 1.130000 0.975000 1.200000 1.055000 ;
      RECT 0.290000 0.905000 1.200000 0.975000 ;
      RECT 0.290000 0.525000 0.360000 0.905000 ;
      RECT 1.130000 0.290000 1.200000 0.905000 ;
      RECT 1.130000 0.220000 1.470000 0.290000 ;
      RECT 1.265000 0.860000 1.335000 0.985000 ;
      RECT 1.265000 0.790000 2.005000 0.860000 ;
      RECT 1.935000 0.860000 2.005000 1.185000 ;
      RECT 1.265000 0.545000 1.335000 0.790000 ;
      RECT 1.265000 0.475000 2.005000 0.545000 ;
      RECT 1.935000 0.185000 2.005000 0.475000 ;
      RECT 2.090000 0.720000 2.160000 1.185000 ;
      RECT 2.090000 0.700000 2.770000 0.720000 ;
      RECT 2.575000 0.720000 2.645000 0.880000 ;
      RECT 1.420000 0.650000 2.770000 0.700000 ;
      RECT 1.420000 0.630000 2.160000 0.650000 ;
      RECT 2.700000 0.350000 2.770000 0.650000 ;
      RECT 2.090000 0.185000 2.160000 0.630000 ;
      RECT 2.630000 0.945000 2.905000 1.015000 ;
      RECT 2.835000 0.440000 2.905000 0.945000 ;
      RECT 2.835000 0.370000 3.270000 0.440000 ;
      RECT 2.835000 0.285000 2.905000 0.370000 ;
      RECT 2.635000 0.215000 2.905000 0.285000 ;
      RECT 2.410000 1.110000 3.040000 1.180000 ;
      RECT 2.970000 0.960000 3.040000 1.110000 ;
      RECT 2.410000 0.785000 2.480000 1.110000 ;
      RECT 2.970000 0.890000 3.400000 0.960000 ;
      RECT 3.330000 0.960000 3.400000 1.185000 ;
      RECT 2.970000 0.575000 3.040000 0.890000 ;
      RECT 2.970000 0.505000 3.405000 0.575000 ;
      RECT 3.335000 0.185000 3.405000 0.505000 ;
      RECT 3.860000 1.030000 3.930000 1.240000 ;
      RECT 3.645000 0.960000 3.930000 1.030000 ;
      RECT 3.645000 0.775000 3.715000 0.960000 ;
      RECT 3.105000 0.640000 3.715000 0.775000 ;
      RECT 3.645000 0.220000 3.715000 0.640000 ;
      RECT 3.645000 0.150000 3.965000 0.220000 ;
      RECT 3.780000 0.490000 3.850000 0.895000 ;
      RECT 3.780000 0.420000 4.050000 0.490000 ;
      RECT 3.980000 0.355000 4.050000 0.420000 ;
      RECT 3.980000 0.285000 4.500000 0.355000 ;
      RECT 4.430000 0.355000 4.500000 1.240000 ;
      RECT 4.430000 0.195000 4.500000 0.285000 ;
  END
END SDFF_X2

MACRO TBUF_X1
  CLASS CORE ;
  FOREIGN TBUF_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.510000 0.495000 0.890000 0.565000 ;
        RECT 0.510000 0.565000 0.580000 0.630000 ;
        RECT 0.820000 0.565000 0.890000 0.730000 ;
    END
    ANTENNAGATEAREA 0.0525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0427 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1768 LAYER metal1 ;
    ANTENNAGATEAREA 0.0525 LAYER metal2 ;
    ANTENNAGATEAREA 0.0525 LAYER metal3 ;
    ANTENNAGATEAREA 0.0525 LAYER metal4 ;
    ANTENNAGATEAREA 0.0525 LAYER metal5 ;
    ANTENNAGATEAREA 0.0525 LAYER metal6 ;
    ANTENNAGATEAREA 0.0525 LAYER metal7 ;
    ANTENNAGATEAREA 0.0525 LAYER metal8 ;
    ANTENNAGATEAREA 0.0525 LAYER metal9 ;
    ANTENNAGATEAREA 0.0525 LAYER metal10 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.200000 0.695000 1.330000 0.920000 ;
    END
    ANTENNAGATEAREA 0.0525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0923 LAYER metal1 ;
    ANTENNAGATEAREA 0.0525 LAYER metal2 ;
    ANTENNAGATEAREA 0.0525 LAYER metal3 ;
    ANTENNAGATEAREA 0.0525 LAYER metal4 ;
    ANTENNAGATEAREA 0.0525 LAYER metal5 ;
    ANTENNAGATEAREA 0.0525 LAYER metal6 ;
    ANTENNAGATEAREA 0.0525 LAYER metal7 ;
    ANTENNAGATEAREA 0.0525 LAYER metal8 ;
    ANTENNAGATEAREA 0.0525 LAYER metal9 ;
    ANTENNAGATEAREA 0.0525 LAYER metal10 ;
  END EN

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.035000 0.425000 0.105000 0.970000 ;
        RECT 0.035000 0.970000 0.140000 1.245000 ;
        RECT 0.035000 0.150000 0.140000 0.425000 ;
    END
    ANTENNADIFFAREA 0.093975 ;
    ANTENNAPARTIALMETALAREA 0.0959 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.520000 1.485000 ;
        RECT 1.190000 1.240000 1.325000 1.315000 ;
        RECT 0.225000 1.145000 0.360000 1.315000 ;
        RECT 0.690000 1.145000 0.760000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.520000 0.085000 ;
        RECT 0.225000 0.085000 0.360000 0.160000 ;
        RECT 0.770000 0.085000 0.905000 0.295000 ;
        RECT 1.150000 0.085000 1.285000 0.295000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.495000 0.905000 0.565000 1.115000 ;
      RECT 0.370000 0.835000 0.565000 0.905000 ;
      RECT 0.370000 0.715000 0.440000 0.835000 ;
      RECT 0.170000 0.645000 0.440000 0.715000 ;
      RECT 0.370000 0.430000 0.440000 0.645000 ;
      RECT 0.370000 0.360000 0.530000 0.430000 ;
      RECT 0.170000 0.495000 0.305000 0.565000 ;
      RECT 0.235000 0.295000 0.305000 0.495000 ;
      RECT 0.235000 0.225000 0.685000 0.295000 ;
      RECT 0.615000 0.295000 0.685000 0.360000 ;
      RECT 0.615000 0.360000 1.135000 0.430000 ;
      RECT 1.065000 0.430000 1.135000 1.040000 ;
      RECT 1.410000 1.175000 1.480000 1.245000 ;
      RECT 0.875000 1.105000 1.480000 1.175000 ;
      RECT 0.875000 1.010000 0.945000 1.105000 ;
      RECT 1.410000 0.435000 1.480000 1.105000 ;
      RECT 0.650000 0.940000 0.945000 1.010000 ;
      RECT 1.345000 0.365000 1.480000 0.435000 ;
      RECT 0.650000 0.645000 0.720000 0.940000 ;
  END
END TBUF_X1

MACRO TBUF_X16
  CLASS CORE ;
  FOREIGN TBUF_X16 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.475000 0.555000 3.740000 0.625000 ;
        RECT 3.670000 0.460000 3.740000 0.555000 ;
        RECT 3.670000 0.390000 4.335000 0.460000 ;
        RECT 4.265000 0.460000 4.335000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3367 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.955000 0.560000 4.120000 0.630000 ;
        RECT 4.050000 0.630000 4.120000 0.725000 ;
        RECT 4.050000 0.725000 4.600000 0.795000 ;
        RECT 4.530000 0.525000 4.600000 0.725000 ;
    END
    ANTENNAGATEAREA 0.15675 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0707 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2808 LAYER metal1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal2 ;
    ANTENNAGATEAREA 0.15675 LAYER metal3 ;
    ANTENNAGATEAREA 0.15675 LAYER metal4 ;
    ANTENNAGATEAREA 0.15675 LAYER metal5 ;
    ANTENNAGATEAREA 0.15675 LAYER metal6 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ;
    ANTENNAGATEAREA 0.15675 LAYER metal8 ;
    ANTENNAGATEAREA 0.15675 LAYER metal9 ;
    ANTENNAGATEAREA 0.15675 LAYER metal10 ;
  END EN

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.240000 0.860000 0.430000 0.930000 ;
        RECT 0.360000 0.700000 0.430000 0.860000 ;
        RECT 0.360000 0.560000 3.030000 0.700000 ;
        RECT 0.620000 0.700000 0.755000 1.005000 ;
        RECT 0.995000 0.700000 1.130000 1.005000 ;
        RECT 1.380000 0.700000 1.515000 1.005000 ;
        RECT 1.755000 0.700000 1.890000 1.005000 ;
        RECT 2.140000 0.700000 2.275000 1.005000 ;
        RECT 2.515000 0.700000 2.650000 1.005000 ;
        RECT 2.895000 0.700000 3.030000 1.005000 ;
        RECT 0.360000 0.430000 0.430000 0.560000 ;
        RECT 0.620000 0.360000 0.755000 0.560000 ;
        RECT 1.000000 0.360000 1.135000 0.560000 ;
        RECT 1.375000 0.360000 1.510000 0.560000 ;
        RECT 1.760000 0.360000 1.895000 0.560000 ;
        RECT 2.135000 0.360000 2.270000 0.560000 ;
        RECT 2.515000 0.360000 2.650000 0.560000 ;
        RECT 2.895000 0.360000 3.030000 0.560000 ;
        RECT 0.240000 0.360000 0.430000 0.430000 ;
    END
    ANTENNADIFFAREA 1.0024 ;
    ANTENNAPARTIALMETALAREA 0.897925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8239 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.940000 1.485000 ;
        RECT 0.050000 1.240000 0.185000 1.315000 ;
        RECT 0.425000 1.240000 0.560000 1.315000 ;
        RECT 0.805000 1.240000 0.940000 1.315000 ;
        RECT 1.185000 1.240000 1.320000 1.315000 ;
        RECT 1.565000 1.240000 1.700000 1.315000 ;
        RECT 1.945000 1.240000 2.080000 1.315000 ;
        RECT 2.325000 1.240000 2.460000 1.315000 ;
        RECT 2.705000 1.240000 2.840000 1.315000 ;
        RECT 3.085000 1.240000 3.220000 1.315000 ;
        RECT 3.465000 1.240000 3.600000 1.315000 ;
        RECT 3.845000 1.240000 3.980000 1.315000 ;
        RECT 4.605000 1.240000 4.740000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.940000 0.085000 ;
        RECT 0.050000 0.085000 0.185000 0.160000 ;
        RECT 0.425000 0.085000 0.560000 0.160000 ;
        RECT 0.805000 0.085000 0.940000 0.160000 ;
        RECT 1.185000 0.085000 1.320000 0.160000 ;
        RECT 1.565000 0.085000 1.700000 0.160000 ;
        RECT 1.945000 0.085000 2.080000 0.160000 ;
        RECT 2.325000 0.085000 2.460000 0.160000 ;
        RECT 2.705000 0.085000 2.840000 0.160000 ;
        RECT 3.085000 0.085000 3.220000 0.160000 ;
        RECT 3.845000 0.085000 3.980000 0.160000 ;
        RECT 4.225000 0.085000 4.360000 0.160000 ;
        RECT 4.605000 0.085000 4.740000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.105000 1.085000 3.790000 1.155000 ;
      RECT 0.105000 0.720000 0.175000 1.085000 ;
      RECT 3.095000 0.430000 3.165000 1.085000 ;
      RECT 0.105000 0.650000 0.295000 0.720000 ;
      RECT 3.095000 0.360000 3.600000 0.430000 ;
      RECT 4.230000 0.860000 4.735000 0.930000 ;
      RECT 4.665000 0.295000 4.735000 0.860000 ;
      RECT 0.105000 0.225000 4.735000 0.295000 ;
      RECT 0.105000 0.295000 0.175000 0.495000 ;
      RECT 0.105000 0.495000 0.290000 0.565000 ;
      RECT 4.825000 1.065000 4.895000 1.250000 ;
      RECT 3.860000 0.995000 4.895000 1.065000 ;
      RECT 3.860000 0.900000 3.930000 0.995000 ;
      RECT 4.825000 0.260000 4.895000 0.995000 ;
      RECT 3.230000 0.830000 3.930000 0.900000 ;
      RECT 3.230000 0.525000 3.300000 0.830000 ;
      RECT 3.805000 0.525000 3.875000 0.830000 ;
  END
END TBUF_X16

MACRO TBUF_X2
  CLASS CORE ;
  FOREIGN TBUF_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.560000 0.965000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.685000 0.285000 1.270000 0.355000 ;
        RECT 1.200000 0.355000 1.270000 0.700000 ;
        RECT 0.685000 0.355000 0.755000 0.660000 ;
        RECT 1.200000 0.700000 1.535000 0.840000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.13335 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4446 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END EN

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.420000 0.130000 0.800000 ;
        RECT 0.060000 0.800000 0.335000 0.870000 ;
        RECT 0.060000 0.350000 0.330000 0.420000 ;
    END
    ANTENNADIFFAREA 0.1253 ;
    ANTENNAPARTIALMETALAREA 0.06475 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2587 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.415000 1.135000 0.485000 1.315000 ;
        RECT 0.975000 1.065000 1.045000 1.315000 ;
        RECT 1.390000 1.065000 1.460000 1.315000 ;
        RECT 0.040000 0.995000 0.110000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.250000 ;
        RECT 0.415000 0.085000 0.485000 0.390000 ;
        RECT 0.910000 0.085000 0.980000 0.200000 ;
        RECT 1.405000 0.085000 1.475000 0.250000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.550000 0.725000 0.705000 0.795000 ;
      RECT 0.550000 0.565000 0.620000 0.725000 ;
      RECT 0.235000 0.495000 0.620000 0.565000 ;
      RECT 0.550000 0.220000 0.620000 0.495000 ;
      RECT 0.550000 0.150000 0.825000 0.220000 ;
      RECT 0.400000 0.925000 1.270000 0.995000 ;
      RECT 0.400000 0.720000 0.470000 0.925000 ;
      RECT 1.065000 0.500000 1.135000 0.925000 ;
      RECT 0.235000 0.650000 0.470000 0.720000 ;
      RECT 1.000000 0.430000 1.135000 0.500000 ;
      RECT 1.600000 0.630000 1.670000 1.250000 ;
      RECT 1.335000 0.560000 1.670000 0.630000 ;
      RECT 1.600000 0.150000 1.670000 0.560000 ;
  END
END TBUF_X2

MACRO TBUF_X4
  CLASS CORE ;
  FOREIGN TBUF_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.350000 0.525000 1.460000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.750000 0.525000 1.840000 0.700000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END EN

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.400000 0.320000 1.065000 ;
        RECT 0.235000 1.065000 0.745000 1.135000 ;
        RECT 0.235000 0.330000 0.745000 0.400000 ;
    END
    ANTENNADIFFAREA 0.2506 ;
    ANTENNAPARTIALMETALAREA 0.127925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4524 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 0.075000 1.205000 0.145000 1.315000 ;
        RECT 0.450000 1.205000 0.520000 1.315000 ;
        RECT 0.830000 1.205000 0.900000 1.315000 ;
        RECT 1.210000 1.205000 1.280000 1.315000 ;
        RECT 1.745000 0.860000 1.815000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.075000 0.085000 0.145000 0.335000 ;
        RECT 0.450000 0.085000 0.520000 0.195000 ;
        RECT 0.830000 0.085000 0.900000 0.195000 ;
        RECT 1.365000 0.085000 1.435000 0.195000 ;
        RECT 1.740000 0.085000 1.810000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.730000 0.725000 1.280000 0.795000 ;
      RECT 0.730000 0.615000 0.800000 0.725000 ;
      RECT 1.210000 0.400000 1.280000 0.725000 ;
      RECT 1.365000 0.965000 1.435000 1.140000 ;
      RECT 0.590000 0.895000 1.630000 0.965000 ;
      RECT 0.590000 0.465000 0.660000 0.895000 ;
      RECT 1.560000 0.400000 1.630000 0.895000 ;
      RECT 0.945000 0.335000 1.015000 0.660000 ;
      RECT 0.945000 0.265000 2.005000 0.335000 ;
      RECT 1.935000 0.335000 2.005000 0.995000 ;
      RECT 1.935000 0.150000 2.005000 0.265000 ;
  END
END TBUF_X4

MACRO TBUF_X8
  CLASS CORE ;
  FOREIGN TBUF_X8 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.42 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.950000 0.560000 2.210000 0.630000 ;
        RECT 2.140000 0.460000 2.210000 0.560000 ;
        RECT 2.140000 0.390000 2.790000 0.460000 ;
        RECT 2.720000 0.460000 2.790000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0847 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3328 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.465000 0.525000 2.600000 0.725000 ;
        RECT 2.465000 0.725000 3.080000 0.795000 ;
        RECT 3.010000 0.525000 3.080000 0.725000 ;
    END
    ANTENNAGATEAREA 0.15675 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08405 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2821 LAYER metal1 ;
    ANTENNAGATEAREA 0.15675 LAYER metal2 ;
    ANTENNAGATEAREA 0.15675 LAYER metal3 ;
    ANTENNAGATEAREA 0.15675 LAYER metal4 ;
    ANTENNAGATEAREA 0.15675 LAYER metal5 ;
    ANTENNAGATEAREA 0.15675 LAYER metal6 ;
    ANTENNAGATEAREA 0.15675 LAYER metal7 ;
    ANTENNAGATEAREA 0.15675 LAYER metal8 ;
    ANTENNAGATEAREA 0.15675 LAYER metal9 ;
    ANTENNAGATEAREA 0.15675 LAYER metal10 ;
  END EN

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.265000 0.775000 1.430000 0.840000 ;
        RECT 0.265000 0.700000 1.425000 0.775000 ;
        RECT 1.360000 0.840000 1.430000 1.010000 ;
        RECT 0.265000 0.840000 0.335000 1.250000 ;
        RECT 0.645000 0.840000 0.715000 1.250000 ;
        RECT 1.020000 0.840000 1.090000 1.250000 ;
        RECT 1.355000 0.445000 1.425000 0.700000 ;
        RECT 0.265000 0.200000 0.335000 0.700000 ;
        RECT 0.645000 0.200000 0.715000 0.700000 ;
        RECT 1.020000 0.200000 1.095000 0.700000 ;
        RECT 1.360000 1.010000 1.505000 1.080000 ;
        RECT 1.355000 0.375000 1.505000 0.445000 ;
    END
    ANTENNADIFFAREA 0.505675 ;
    ANTENNAPARTIALMETALAREA 0.406725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2363 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.420000 1.485000 ;
        RECT 2.320000 1.150000 2.455000 1.315000 ;
        RECT 3.085000 1.130000 3.220000 1.315000 ;
        RECT 0.415000 1.010000 0.550000 1.315000 ;
        RECT 1.590000 0.995000 1.660000 1.315000 ;
        RECT 1.970000 0.995000 2.040000 1.315000 ;
        RECT 0.070000 0.975000 0.140000 1.315000 ;
        RECT 0.830000 0.975000 0.900000 1.315000 ;
        RECT 1.210000 0.975000 1.280000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.420000 0.085000 ;
        RECT 0.070000 0.085000 0.140000 0.410000 ;
        RECT 0.415000 0.085000 0.550000 0.375000 ;
        RECT 0.800000 0.085000 0.935000 0.160000 ;
        RECT 1.180000 0.085000 1.315000 0.160000 ;
        RECT 1.560000 0.085000 1.695000 0.160000 ;
        RECT 2.320000 0.085000 2.455000 0.160000 ;
        RECT 2.700000 0.085000 2.835000 0.160000 ;
        RECT 3.090000 0.085000 3.225000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.780000 0.930000 1.850000 1.250000 ;
      RECT 1.570000 0.860000 2.230000 0.930000 ;
      RECT 2.160000 0.930000 2.230000 1.250000 ;
      RECT 1.570000 0.750000 1.640000 0.860000 ;
      RECT 1.490000 0.615000 1.640000 0.750000 ;
      RECT 1.570000 0.460000 1.640000 0.615000 ;
      RECT 1.570000 0.390000 2.075000 0.460000 ;
      RECT 2.705000 0.860000 3.215000 0.930000 ;
      RECT 3.145000 0.295000 3.215000 0.860000 ;
      RECT 1.205000 0.225000 3.215000 0.295000 ;
      RECT 1.205000 0.295000 1.275000 0.600000 ;
      RECT 3.305000 1.065000 3.375000 1.250000 ;
      RECT 2.295000 0.995000 3.375000 1.065000 ;
      RECT 2.295000 0.795000 2.365000 0.995000 ;
      RECT 3.305000 0.200000 3.375000 0.995000 ;
      RECT 1.705000 0.725000 2.365000 0.795000 ;
      RECT 1.705000 0.525000 1.775000 0.725000 ;
      RECT 2.275000 0.525000 2.365000 0.725000 ;
  END
END TBUF_X8

MACRO TINV_X1
  CLASS CORE ;
  FOREIGN TINV_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.175000 0.625000 0.245000 0.840000 ;
        RECT 0.175000 0.840000 0.520000 0.980000 ;
        RECT 0.450000 0.720000 0.520000 0.840000 ;
        RECT 0.450000 0.650000 0.585000 0.720000 ;
    END
    ANTENNAGATEAREA 0.05325 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0812 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2483 LAYER metal1 ;
    ANTENNAGATEAREA 0.05325 LAYER metal2 ;
    ANTENNAGATEAREA 0.05325 LAYER metal3 ;
    ANTENNAGATEAREA 0.05325 LAYER metal4 ;
    ANTENNAGATEAREA 0.05325 LAYER metal5 ;
    ANTENNAGATEAREA 0.05325 LAYER metal6 ;
    ANTENNAGATEAREA 0.05325 LAYER metal7 ;
    ANTENNAGATEAREA 0.05325 LAYER metal8 ;
    ANTENNAGATEAREA 0.05325 LAYER metal9 ;
    ANTENNAGATEAREA 0.05325 LAYER metal10 ;
  END EN

  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.420000 0.380000 0.560000 ;
        RECT 0.310000 0.560000 0.380000 0.600000 ;
    END
    ANTENNAGATEAREA 0.04475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.04475 LAYER metal2 ;
    ANTENNAGATEAREA 0.04475 LAYER metal3 ;
    ANTENNAGATEAREA 0.04475 LAYER metal4 ;
    ANTENNAGATEAREA 0.04475 LAYER metal5 ;
    ANTENNAGATEAREA 0.04475 LAYER metal6 ;
    ANTENNAGATEAREA 0.04475 LAYER metal7 ;
    ANTENNAGATEAREA 0.04475 LAYER metal8 ;
    ANTENNAGATEAREA 0.04475 LAYER metal9 ;
    ANTENNAGATEAREA 0.04475 LAYER metal10 ;
  END I

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.840000 0.720000 1.240000 ;
        RECT 0.650000 0.155000 0.720000 0.840000 ;
    END
    ANTENNADIFFAREA 0.093975 ;
    ANTENNAPARTIALMETALAREA 0.08395 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3055 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.225000 1.065000 0.295000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.450000 0.495000 0.585000 0.565000 ;
      RECT 0.450000 0.345000 0.520000 0.495000 ;
      RECT 0.040000 0.275000 0.520000 0.345000 ;
      RECT 0.040000 0.345000 0.110000 1.240000 ;
      RECT 0.040000 0.195000 0.110000 0.275000 ;
  END
END TINV_X1

MACRO TLAT_X1
  CLASS CORE ;
  FOREIGN TLAT_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.585000 0.730000 0.840000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0255 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0923 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185000 0.745000 0.320000 0.980000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.031725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0962 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END G

  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.815000 0.500000 2.275000 0.570000 ;
        RECT 1.815000 0.570000 2.030000 0.700000 ;
    END
    ANTENNAGATEAREA 0.044 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.06015 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1716 LAYER metal1 ;
    ANTENNAGATEAREA 0.044 LAYER metal2 ;
    ANTENNAGATEAREA 0.044 LAYER metal3 ;
    ANTENNAGATEAREA 0.044 LAYER metal4 ;
    ANTENNAGATEAREA 0.044 LAYER metal5 ;
    ANTENNAGATEAREA 0.044 LAYER metal6 ;
    ANTENNAGATEAREA 0.044 LAYER metal7 ;
    ANTENNAGATEAREA 0.044 LAYER metal8 ;
    ANTENNAGATEAREA 0.044 LAYER metal9 ;
    ANTENNAGATEAREA 0.044 LAYER metal10 ;
  END OE

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.265000 1.010000 2.410000 1.215000 ;
        RECT 2.340000 0.425000 2.410000 1.010000 ;
        RECT 2.265000 0.220000 2.410000 0.425000 ;
    END
    ANTENNADIFFAREA 0.111875 ;
    ANTENNAPARTIALMETALAREA 0.1004 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3159 LAYER metal1 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 1.305000 1.080000 1.440000 1.315000 ;
        RECT 0.235000 1.045000 0.305000 1.315000 ;
        RECT 0.585000 1.040000 0.655000 1.315000 ;
        RECT 1.870000 0.975000 1.940000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.235000 0.085000 0.305000 0.320000 ;
        RECT 0.585000 0.085000 0.655000 0.460000 ;
        RECT 1.335000 0.085000 1.405000 0.320000 ;
        RECT 1.870000 0.085000 1.940000 0.320000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.050000 0.595000 0.120000 1.250000 ;
      RECT 0.050000 0.460000 0.365000 0.595000 ;
      RECT 0.050000 0.185000 0.120000 0.460000 ;
      RECT 0.430000 0.975000 0.500000 1.250000 ;
      RECT 0.430000 0.905000 0.945000 0.975000 ;
      RECT 0.875000 0.510000 0.945000 0.905000 ;
      RECT 0.430000 0.185000 0.500000 0.905000 ;
      RECT 0.930000 1.070000 1.090000 1.140000 ;
      RECT 1.020000 0.880000 1.090000 1.070000 ;
      RECT 1.020000 0.745000 1.465000 0.880000 ;
      RECT 1.020000 0.290000 1.090000 0.745000 ;
      RECT 0.930000 0.220000 1.090000 0.290000 ;
      RECT 1.530000 0.650000 1.600000 1.185000 ;
      RECT 1.260000 0.515000 1.600000 0.650000 ;
      RECT 1.530000 0.185000 1.600000 0.515000 ;
      RECT 1.680000 0.855000 1.750000 1.245000 ;
      RECT 1.680000 0.775000 2.275000 0.855000 ;
      RECT 2.140000 0.650000 2.275000 0.775000 ;
      RECT 1.680000 0.185000 1.750000 0.775000 ;
  END
END TLAT_X1

MACRO NAND4_X1
  CLASS CORE ;
  FOREIGN NAND4_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.420000 0.555000 0.660000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0276 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0923 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.420000 0.375000 0.660000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.03 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0949 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.420000 0.185000 0.660000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.03 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0949 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.840000 0.700000 0.910000 ;
        RECT 0.235000 0.910000 0.305000 1.250000 ;
        RECT 0.615000 0.910000 0.700000 1.250000 ;
        RECT 0.630000 0.425000 0.700000 0.840000 ;
        RECT 0.630000 0.355000 0.865000 0.425000 ;
        RECT 0.795000 0.150000 0.865000 0.355000 ;
    END
    ANTENNADIFFAREA 0.219975 ;
    ANTENNAPARTIALMETALAREA 0.1451 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5382 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.355000 ;
    END
  END VSS
END NAND4_X1

MACRO NAND4_X2
  CLASS CORE ;
  FOREIGN NAND4_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.810000 0.420000 0.945000 0.625000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.027675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0884 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.285000 1.270000 0.355000 ;
        RECT 0.575000 0.355000 0.645000 0.660000 ;
        RECT 1.145000 0.355000 1.270000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.108125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3575 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.390000 0.525000 0.510000 0.725000 ;
        RECT 0.390000 0.725000 1.405000 0.795000 ;
        RECT 1.335000 0.525000 1.405000 0.725000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.10905 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3861 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.320000 0.860000 ;
        RECT 0.195000 0.860000 1.590000 0.930000 ;
        RECT 1.520000 0.525000 1.590000 0.860000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.162975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5551 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.995000 1.510000 1.065000 ;
        RECT 0.060000 0.460000 0.130000 0.995000 ;
        RECT 0.235000 1.065000 0.370000 1.250000 ;
        RECT 0.615000 1.065000 0.750000 1.250000 ;
        RECT 0.995000 1.065000 1.130000 1.250000 ;
        RECT 1.375000 1.065000 1.510000 1.250000 ;
        RECT 0.060000 0.390000 0.355000 0.460000 ;
        RECT 0.285000 0.220000 0.355000 0.390000 ;
        RECT 0.285000 0.150000 0.940000 0.220000 ;
    END
    ANTENNADIFFAREA 0.4109 ;
    ANTENNAPARTIALMETALAREA 0.31725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.0179 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.080000 1.130000 0.150000 1.315000 ;
        RECT 0.455000 1.130000 0.525000 1.315000 ;
        RECT 0.835000 1.130000 0.905000 1.315000 ;
        RECT 1.215000 1.130000 1.285000 1.315000 ;
        RECT 1.595000 1.065000 1.665000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.250000 ;
        RECT 1.595000 0.085000 1.665000 0.390000 ;
    END
  END VSS
END NAND4_X2

MACRO NAND4_X4
  CLASS CORE ;
  FOREIGN NAND4_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.42 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.405000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.018375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.170000 0.525000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.150000 0.525000 2.220000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.910000 0.525000 2.980000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.090000 0.840000 3.340000 0.980000 ;
        RECT 0.090000 0.980000 0.160000 1.155000 ;
        RECT 0.460000 0.980000 0.530000 1.155000 ;
        RECT 0.840000 0.980000 0.910000 1.155000 ;
        RECT 1.220000 0.980000 1.290000 1.155000 ;
        RECT 1.680000 0.980000 1.750000 1.155000 ;
        RECT 2.130000 0.980000 2.200000 1.155000 ;
        RECT 2.510000 0.980000 2.580000 1.155000 ;
        RECT 2.890000 0.980000 2.960000 1.155000 ;
        RECT 3.270000 0.980000 3.340000 1.155000 ;
        RECT 0.685000 0.355000 0.755000 0.840000 ;
        RECT 0.225000 0.285000 0.755000 0.355000 ;
    END
    ANTENNADIFFAREA 0.9604 ;
    ANTENNAPARTIALMETALAREA 0.6363 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5548 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.420000 1.485000 ;
        RECT 0.240000 1.095000 0.375000 1.315000 ;
        RECT 0.620000 1.095000 0.755000 1.315000 ;
        RECT 1.000000 1.095000 1.135000 1.315000 ;
        RECT 1.380000 1.095000 1.515000 1.315000 ;
        RECT 1.910000 1.095000 2.045000 1.315000 ;
        RECT 2.290000 1.095000 2.425000 1.315000 ;
        RECT 2.670000 1.095000 2.805000 1.315000 ;
        RECT 3.050000 1.095000 3.185000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.420000 0.085000 ;
        RECT 2.670000 0.085000 2.805000 0.300000 ;
        RECT 3.050000 0.085000 3.185000 0.300000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.090000 0.220000 0.160000 0.460000 ;
      RECT 0.090000 0.150000 1.670000 0.220000 ;
      RECT 0.840000 0.220000 0.910000 0.460000 ;
      RECT 1.600000 0.220000 1.670000 0.460000 ;
      RECT 1.380000 0.525000 2.045000 0.595000 ;
      RECT 1.380000 0.355000 1.515000 0.525000 ;
      RECT 1.910000 0.355000 2.045000 0.525000 ;
      RECT 1.005000 0.285000 1.515000 0.355000 ;
      RECT 1.910000 0.285000 2.425000 0.355000 ;
      RECT 1.760000 0.220000 1.830000 0.460000 ;
      RECT 1.760000 0.150000 2.580000 0.220000 ;
      RECT 2.510000 0.220000 2.580000 0.390000 ;
      RECT 2.510000 0.390000 3.340000 0.460000 ;
      RECT 2.890000 0.185000 2.960000 0.390000 ;
      RECT 3.270000 0.185000 3.340000 0.390000 ;
  END
END NAND4_X4

MACRO NOR2_X1
  CLASS CORE ;
  FOREIGN NOR2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.150000 0.320000 0.975000 ;
        RECT 0.250000 0.975000 0.500000 1.045000 ;
        RECT 0.430000 1.045000 0.500000 1.250000 ;
    END
    ANTENNADIFFAREA 0.12425 ;
    ANTENNAPARTIALMETALAREA 0.0896 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.570000 1.485000 ;
        RECT 0.055000 0.975000 0.125000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.570000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.425000 ;
        RECT 0.430000 0.085000 0.500000 0.425000 ;
    END
  END VSS
END NOR2_X1

MACRO NOR2_X2
  CLASS CORE ;
  FOREIGN NOR2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.420000 0.510000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.265000 0.725000 ;
        RECT 0.195000 0.725000 0.890000 0.795000 ;
        RECT 0.760000 0.525000 0.890000 0.725000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08865 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3029 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.260000 0.750000 0.330000 ;
        RECT 0.060000 0.330000 0.130000 0.910000 ;
        RECT 0.060000 0.910000 0.525000 0.980000 ;
        RECT 0.455000 0.980000 0.525000 1.250000 ;
    END
    ANTENNADIFFAREA 0.2044 ;
    ANTENNAPARTIALMETALAREA 0.14035 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5395 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.080000 1.045000 0.150000 1.315000 ;
        RECT 0.835000 1.045000 0.905000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.195000 ;
        RECT 0.455000 0.085000 0.525000 0.195000 ;
        RECT 0.835000 0.085000 0.905000 0.335000 ;
    END
  END VSS
END NOR2_X2

MACRO NOR2_X4
  CLASS CORE ;
  FOREIGN NOR2_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.590000 0.420000 1.160000 0.490000 ;
        RECT 0.590000 0.490000 0.700000 0.660000 ;
        RECT 1.090000 0.490000 1.160000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0705 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2548 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.215000 0.525000 0.285000 0.910000 ;
        RECT 0.215000 0.910000 1.535000 0.980000 ;
        RECT 0.805000 0.560000 0.940000 0.910000 ;
        RECT 1.465000 0.525000 1.535000 0.910000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.19355 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6526 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.240000 0.280000 1.510000 0.350000 ;
        RECT 0.440000 0.350000 0.525000 0.845000 ;
        RECT 1.225000 0.350000 1.295000 0.845000 ;
    END
    ANTENNADIFFAREA 0.4088 ;
    ANTENNAPARTIALMETALAREA 0.165625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6058 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.835000 1.045000 0.905000 1.315000 ;
        RECT 0.080000 0.710000 0.150000 1.315000 ;
        RECT 1.600000 0.710000 1.670000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.390000 ;
        RECT 0.455000 0.085000 0.525000 0.195000 ;
        RECT 0.835000 0.085000 0.905000 0.195000 ;
        RECT 1.215000 0.085000 1.285000 0.195000 ;
        RECT 1.595000 0.085000 1.665000 0.390000 ;
    END
  END VSS
END NOR2_X4

MACRO NOR3_X1
  CLASS CORE ;
  FOREIGN NOR3_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.545000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.018375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.175000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.020125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0754 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.150000 0.305000 0.355000 ;
        RECT 0.235000 0.355000 0.700000 0.425000 ;
        RECT 0.610000 0.425000 0.700000 1.000000 ;
        RECT 0.610000 0.150000 0.700000 0.355000 ;
    END
    ANTENNADIFFAREA 0.167825 ;
    ANTENNAPARTIALMETALAREA 0.1171 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3952 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.220000 ;
    END
  END VSS
END NOR3_X1

MACRO NOR3_X2
  CLASS CORE ;
  FOREIGN NOR3_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.620000 0.560000 0.755000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.390000 0.425000 0.990000 0.495000 ;
        RECT 0.390000 0.495000 0.510000 0.700000 ;
        RECT 0.920000 0.495000 0.990000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.07815 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2704 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.265000 0.770000 ;
        RECT 0.195000 0.770000 1.270000 0.840000 ;
        RECT 1.145000 0.525000 1.270000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.123025 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4251 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.285000 1.130000 0.355000 ;
        RECT 0.060000 0.355000 0.130000 0.905000 ;
        RECT 0.060000 0.905000 0.715000 0.975000 ;
        RECT 0.645000 0.975000 0.715000 1.180000 ;
    END
    ANTENNADIFFAREA 0.2625 ;
    ANTENNAPARTIALMETALAREA 0.1736 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.663 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.080000 1.065000 0.150000 1.315000 ;
        RECT 1.215000 1.065000 1.285000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.195000 ;
        RECT 0.455000 0.085000 0.525000 0.195000 ;
        RECT 0.835000 0.085000 0.905000 0.195000 ;
        RECT 1.215000 0.085000 1.285000 0.335000 ;
    END
  END VSS
END NOR3_X2

MACRO NOR3_X4
  CLASS CORE ;
  FOREIGN NOR3_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.185000 0.525000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.130000 0.525000 2.230000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.150000 0.305000 0.390000 ;
        RECT 0.235000 0.390000 2.380000 0.460000 ;
        RECT 0.235000 0.460000 0.320000 0.765000 ;
        RECT 0.605000 0.150000 0.675000 0.390000 ;
        RECT 0.985000 0.150000 1.055000 0.390000 ;
        RECT 1.365000 0.150000 1.435000 0.390000 ;
        RECT 1.930000 0.150000 2.000000 0.390000 ;
        RECT 2.310000 0.150000 2.380000 0.390000 ;
        RECT 0.235000 0.765000 0.675000 0.835000 ;
        RECT 0.235000 0.835000 0.305000 1.115000 ;
        RECT 0.605000 0.835000 0.675000 1.115000 ;
    END
    ANTENNADIFFAREA 0.525 ;
    ANTENNAPARTIALMETALAREA 0.346875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2857 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.660000 1.485000 ;
        RECT 2.090000 0.935000 2.225000 1.315000 ;
        RECT 1.745000 0.900000 1.815000 1.315000 ;
        RECT 2.500000 0.900000 2.570000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.660000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.385000 0.085000 0.520000 0.325000 ;
        RECT 0.765000 0.085000 0.900000 0.325000 ;
        RECT 1.145000 0.085000 1.280000 0.325000 ;
        RECT 1.525000 0.085000 1.850000 0.325000 ;
        RECT 2.090000 0.085000 2.225000 0.325000 ;
        RECT 2.505000 0.085000 2.575000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 1.180000 1.625000 1.250000 ;
      RECT 0.045000 0.900000 0.115000 1.180000 ;
      RECT 0.415000 0.900000 0.485000 1.180000 ;
      RECT 0.795000 0.900000 0.865000 1.180000 ;
      RECT 1.175000 0.900000 1.245000 1.180000 ;
      RECT 1.555000 0.900000 1.625000 1.180000 ;
      RECT 0.995000 0.835000 1.065000 1.115000 ;
      RECT 0.995000 0.765000 2.380000 0.835000 ;
      RECT 1.365000 0.835000 1.435000 1.115000 ;
      RECT 1.930000 0.835000 2.000000 1.175000 ;
      RECT 2.310000 0.835000 2.380000 1.175000 ;
  END
END NOR3_X4

MACRO NOR4_X1
  CLASS CORE ;
  FOREIGN NOR4_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.150000 0.305000 0.355000 ;
        RECT 0.235000 0.355000 0.700000 0.425000 ;
        RECT 0.630000 0.425000 0.700000 0.975000 ;
        RECT 0.610000 0.150000 0.700000 0.355000 ;
        RECT 0.630000 0.975000 0.865000 1.045000 ;
        RECT 0.795000 1.045000 0.865000 1.250000 ;
    END
    ANTENNADIFFAREA 0.18235 ;
    ANTENNAPARTIALMETALAREA 0.13465 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5031 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.425000 ;
    END
  END VSS
END NOR4_X1

MACRO NOR4_X2
  CLASS CORE ;
  FOREIGN NOR4_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.810000 0.560000 0.945000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.570000 0.420000 1.180000 0.490000 ;
        RECT 0.570000 0.490000 0.700000 0.700000 ;
        RECT 1.110000 0.490000 1.180000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0819 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2756 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.380000 0.525000 0.450000 0.765000 ;
        RECT 0.380000 0.765000 1.460000 0.835000 ;
        RECT 1.330000 0.525000 1.460000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1236 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4238 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.200000 0.525000 0.270000 0.910000 ;
        RECT 0.200000 0.910000 1.650000 0.980000 ;
        RECT 1.525000 0.840000 1.650000 0.910000 ;
        RECT 1.525000 0.525000 1.595000 0.840000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.15925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5954 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.055000 0.260000 1.475000 0.330000 ;
        RECT 0.055000 0.330000 0.130000 1.055000 ;
        RECT 1.405000 0.330000 1.475000 0.425000 ;
        RECT 1.405000 0.150000 1.475000 0.260000 ;
        RECT 0.055000 1.055000 0.940000 1.125000 ;
    END
    ANTENNADIFFAREA 0.3206 ;
    ANTENNAPARTIALMETALAREA 0.230075 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.858 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.080000 1.205000 0.150000 1.315000 ;
        RECT 1.595000 1.065000 1.665000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.195000 ;
        RECT 0.425000 0.085000 0.560000 0.160000 ;
        RECT 0.805000 0.085000 0.940000 0.160000 ;
        RECT 1.185000 0.085000 1.320000 0.160000 ;
        RECT 1.595000 0.085000 1.665000 0.335000 ;
    END
  END VSS
END NOR4_X2

MACRO NOR4_X4
  CLASS CORE ;
  FOREIGN NOR4_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.42 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.180000 0.525000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.150000 0.525000 2.245000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.016625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.910000 0.525000 3.000000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.150000 0.305000 0.390000 ;
        RECT 0.235000 0.390000 3.375000 0.460000 ;
        RECT 0.235000 0.460000 0.320000 0.765000 ;
        RECT 0.605000 0.150000 0.675000 0.390000 ;
        RECT 0.985000 0.150000 1.055000 0.390000 ;
        RECT 1.370000 0.150000 1.440000 0.390000 ;
        RECT 1.790000 0.150000 1.860000 0.390000 ;
        RECT 2.165000 0.150000 2.235000 0.390000 ;
        RECT 2.545000 0.150000 2.615000 0.390000 ;
        RECT 2.925000 0.150000 2.995000 0.390000 ;
        RECT 3.305000 0.150000 3.375000 0.390000 ;
        RECT 0.235000 0.765000 0.675000 0.835000 ;
        RECT 0.235000 0.835000 0.305000 1.115000 ;
        RECT 0.605000 0.835000 0.675000 1.115000 ;
    END
    ANTENNADIFFAREA 0.67025 ;
    ANTENNAPARTIALMETALAREA 0.466925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7316 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.420000 1.485000 ;
        RECT 2.705000 0.935000 2.840000 1.315000 ;
        RECT 3.085000 0.935000 3.220000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.420000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.360000 ;
        RECT 0.385000 0.085000 0.520000 0.325000 ;
        RECT 0.765000 0.085000 0.900000 0.325000 ;
        RECT 1.145000 0.085000 1.280000 0.325000 ;
        RECT 1.525000 0.085000 1.660000 0.325000 ;
        RECT 1.945000 0.085000 2.080000 0.325000 ;
        RECT 2.325000 0.085000 2.460000 0.325000 ;
        RECT 2.705000 0.085000 2.840000 0.325000 ;
        RECT 3.085000 0.085000 3.220000 0.325000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 1.180000 0.865000 1.250000 ;
      RECT 0.045000 0.900000 0.115000 1.180000 ;
      RECT 0.415000 0.900000 0.485000 1.180000 ;
      RECT 0.795000 0.835000 0.865000 1.180000 ;
      RECT 0.795000 0.765000 1.625000 0.835000 ;
      RECT 1.175000 0.835000 1.245000 1.115000 ;
      RECT 1.555000 0.835000 1.625000 1.115000 ;
      RECT 0.995000 1.180000 2.425000 1.250000 ;
      RECT 0.995000 0.900000 1.065000 1.180000 ;
      RECT 1.365000 0.900000 1.435000 1.180000 ;
      RECT 1.975000 0.900000 2.045000 1.180000 ;
      RECT 2.355000 0.900000 2.425000 1.180000 ;
      RECT 1.795000 0.835000 1.865000 1.115000 ;
      RECT 1.795000 0.765000 3.375000 0.835000 ;
      RECT 2.165000 0.835000 2.235000 1.115000 ;
      RECT 2.545000 0.835000 2.615000 1.175000 ;
      RECT 2.925000 0.835000 2.995000 1.175000 ;
      RECT 3.305000 0.835000 3.375000 1.175000 ;
  END
END NOR4_X4

MACRO OAI211_X1
  CLASS CORE ;
  FOREIGN OAI211_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.790000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.400000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.285000 0.335000 0.780000 ;
        RECT 0.250000 0.780000 0.905000 0.850000 ;
        RECT 0.250000 0.850000 0.525000 0.855000 ;
        RECT 0.835000 0.850000 0.905000 1.055000 ;
        RECT 0.455000 0.855000 0.525000 1.055000 ;
    END
    ANTENNADIFFAREA 0.21245 ;
    ANTENNAPARTIALMETALAREA 0.11765 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4238 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.080000 1.040000 0.150000 1.315000 ;
        RECT 0.645000 1.040000 0.715000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.835000 0.085000 0.905000 0.460000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085000 0.220000 0.155000 0.425000 ;
      RECT 0.085000 0.150000 0.525000 0.220000 ;
      RECT 0.455000 0.220000 0.525000 0.425000 ;
  END
END OAI211_X1

MACRO OAI211_X2
  CLASS CORE ;
  FOREIGN OAI211_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.185000 0.525000 0.320000 0.765000 ;
        RECT 0.185000 0.765000 0.755000 0.835000 ;
        RECT 0.685000 0.525000 0.755000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0891 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2912 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.530000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.190000 0.525000 1.290000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.960000 0.525000 1.030000 0.770000 ;
        RECT 0.960000 0.770000 1.650000 0.840000 ;
        RECT 1.525000 0.525000 1.650000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.096075 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.270000 0.905000 1.285000 0.975000 ;
        RECT 0.270000 0.975000 0.340000 1.250000 ;
        RECT 0.645000 0.975000 0.715000 1.250000 ;
        RECT 1.215000 0.975000 1.285000 1.250000 ;
        RECT 0.820000 0.460000 0.890000 0.905000 ;
        RECT 0.820000 0.390000 1.510000 0.460000 ;
    END
    ANTENNADIFFAREA 0.38395 ;
    ANTENNAPARTIALMETALAREA 0.20825 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7917 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.080000 1.040000 0.150000 1.315000 ;
        RECT 0.455000 1.040000 0.525000 1.315000 ;
        RECT 0.835000 1.040000 0.905000 1.315000 ;
        RECT 1.595000 1.040000 1.665000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.450000 0.085000 0.520000 0.320000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.080000 0.390000 0.660000 0.460000 ;
      RECT 0.590000 0.255000 0.660000 0.390000 ;
      RECT 0.080000 0.185000 0.150000 0.390000 ;
      RECT 0.590000 0.185000 1.665000 0.255000 ;
      RECT 1.595000 0.255000 1.665000 0.460000 ;
  END
END OAI211_X2

MACRO OAI211_X4
  CLASS CORE ;
  FOREIGN OAI211_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.125000 0.390000 1.520000 0.460000 ;
        RECT 0.125000 0.460000 0.195000 0.660000 ;
        RECT 0.805000 0.460000 0.875000 0.660000 ;
        RECT 1.390000 0.460000 1.520000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.15165 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5369 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.420000 0.525000 0.510000 0.770000 ;
        RECT 0.420000 0.770000 1.245000 0.840000 ;
        RECT 1.175000 0.525000 1.245000 0.770000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09695 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3601 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.910000 0.560000 2.045000 0.770000 ;
        RECT 1.910000 0.770000 2.800000 0.840000 ;
        RECT 2.665000 0.560000 2.800000 0.770000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.119 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3588 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.670000 0.425000 3.035000 0.495000 ;
        RECT 1.670000 0.495000 1.740000 0.660000 ;
        RECT 2.310000 0.495000 2.410000 0.700000 ;
        RECT 2.965000 0.495000 3.035000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.13915 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5122 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.905000 3.170000 0.975000 ;
        RECT 0.235000 0.975000 0.305000 1.250000 ;
        RECT 0.605000 0.975000 0.675000 1.250000 ;
        RECT 0.985000 0.975000 1.055000 1.250000 ;
        RECT 1.365000 0.975000 1.435000 1.250000 ;
        RECT 1.935000 0.975000 2.005000 1.250000 ;
        RECT 2.695000 0.975000 2.765000 1.250000 ;
        RECT 3.100000 0.360000 3.170000 0.905000 ;
        RECT 1.720000 0.290000 3.170000 0.360000 ;
    END
    ANTENNADIFFAREA 0.7616 ;
    ANTENNAPARTIALMETALAREA 0.4606 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.729 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.230000 1.485000 ;
        RECT 0.040000 1.040000 0.110000 1.315000 ;
        RECT 0.415000 1.040000 0.485000 1.315000 ;
        RECT 0.795000 1.040000 0.865000 1.315000 ;
        RECT 1.175000 1.040000 1.245000 1.315000 ;
        RECT 1.555000 1.040000 1.625000 1.315000 ;
        RECT 2.315000 1.040000 2.385000 1.315000 ;
        RECT 3.075000 1.040000 3.145000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.230000 0.085000 ;
        RECT 0.385000 0.085000 0.520000 0.160000 ;
        RECT 1.145000 0.085000 1.280000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.225000 1.625000 0.295000 ;
      RECT 1.555000 0.220000 1.625000 0.225000 ;
      RECT 0.045000 0.150000 0.115000 0.225000 ;
      RECT 1.555000 0.150000 3.180000 0.220000 ;
  END
END OAI211_X4

MACRO OAI21_X1
  CLASS CORE ;
  FOREIGN OAI21_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.285000 0.320000 0.765000 ;
        RECT 0.250000 0.765000 0.510000 0.835000 ;
        RECT 0.440000 0.835000 0.510000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.08085 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3185 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.065000 0.975000 0.135000 1.315000 ;
        RECT 0.630000 0.975000 0.700000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.630000 0.085000 0.700000 0.460000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.070000 0.220000 0.140000 0.425000 ;
      RECT 0.070000 0.150000 0.510000 0.220000 ;
      RECT 0.440000 0.220000 0.510000 0.425000 ;
  END
END OAI21_X1

MACRO OAI21_X2
  CLASS CORE ;
  FOREIGN OAI21_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.190000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.570000 0.770000 ;
        RECT 0.440000 0.770000 1.135000 0.840000 ;
        RECT 1.065000 0.525000 1.135000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09765 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3263 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.905000 1.270000 0.975000 ;
        RECT 0.235000 0.975000 0.305000 1.250000 ;
        RECT 0.795000 0.975000 0.865000 1.250000 ;
        RECT 1.200000 0.425000 1.270000 0.905000 ;
        RECT 0.580000 0.355000 1.270000 0.425000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.19285 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7345 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.040000 1.040000 0.110000 1.315000 ;
        RECT 0.415000 1.040000 0.485000 1.315000 ;
        RECT 1.175000 1.040000 1.245000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.355000 0.485000 0.425000 ;
      RECT 0.415000 0.220000 0.485000 0.355000 ;
      RECT 0.045000 0.150000 0.115000 0.355000 ;
      RECT 0.415000 0.150000 1.280000 0.220000 ;
  END
END OAI21_X2

MACRO OAI21_X4
  CLASS CORE ;
  FOREIGN OAI21_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.430000 0.525000 0.515000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.150000 0.560000 1.285000 0.690000 ;
        RECT 1.150000 0.690000 2.040000 0.760000 ;
        RECT 1.905000 0.560000 2.040000 0.690000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0974 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3172 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.910000 0.420000 2.275000 0.490000 ;
        RECT 0.910000 0.490000 0.980000 0.660000 ;
        RECT 1.525000 0.490000 1.660000 0.625000 ;
        RECT 2.150000 0.490000 2.275000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.146925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4966 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.845000 2.410000 0.915000 ;
        RECT 0.235000 0.915000 0.305000 1.190000 ;
        RECT 0.605000 0.915000 0.675000 1.190000 ;
        RECT 1.175000 0.915000 1.245000 1.190000 ;
        RECT 1.935000 0.915000 2.005000 1.190000 ;
        RECT 2.340000 0.355000 2.410000 0.845000 ;
        RECT 0.960000 0.285000 2.410000 0.355000 ;
    END
    ANTENNADIFFAREA 0.5852 ;
    ANTENNAPARTIALMETALAREA 0.36505 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3741 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.040000 1.040000 0.110000 1.315000 ;
        RECT 0.415000 1.040000 0.485000 1.315000 ;
        RECT 0.795000 1.040000 0.865000 1.315000 ;
        RECT 1.555000 1.040000 1.625000 1.315000 ;
        RECT 2.315000 1.040000 2.385000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.355000 0.830000 0.425000 ;
      RECT 0.760000 0.220000 0.830000 0.355000 ;
      RECT 0.045000 0.150000 0.115000 0.355000 ;
      RECT 0.420000 0.150000 0.490000 0.355000 ;
      RECT 0.760000 0.150000 2.420000 0.220000 ;
  END
END OAI21_X4

MACRO OAI221_X1
  CLASS CORE ;
  FOREIGN OAI221_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.740000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.850000 1.055000 0.920000 ;
        RECT 0.425000 0.920000 0.495000 1.250000 ;
        RECT 0.985000 0.920000 1.055000 1.250000 ;
        RECT 0.805000 0.400000 0.890000 0.850000 ;
    END
    ANTENNADIFFAREA 0.21245 ;
    ANTENNAPARTIALMETALAREA 0.12855 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4706 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.040000 1.040000 0.110000 1.315000 ;
        RECT 0.605000 1.040000 0.675000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.355000 0.485000 0.425000 ;
      RECT 0.045000 0.150000 0.115000 0.355000 ;
      RECT 0.415000 0.150000 0.485000 0.355000 ;
      RECT 0.615000 0.220000 0.685000 0.425000 ;
      RECT 0.615000 0.150000 1.055000 0.220000 ;
      RECT 0.985000 0.220000 1.055000 0.425000 ;
  END
END OAI221_X1

MACRO OAI221_X2
  CLASS CORE ;
  FOREIGN OAI221_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955000 0.525000 1.025000 0.900000 ;
        RECT 0.955000 0.900000 2.030000 0.970000 ;
        RECT 1.930000 0.525000 2.030000 0.900000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.139 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4927 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.155000 0.525000 1.225000 0.765000 ;
        RECT 1.155000 0.765000 1.840000 0.835000 ;
        RECT 1.715000 0.525000 1.840000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09475 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3211 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.380000 0.525000 1.480000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.525000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.265000 0.770000 ;
        RECT 0.195000 0.770000 0.890000 0.840000 ;
        RECT 0.760000 0.525000 0.890000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09765 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3263 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 1.035000 1.890000 1.105000 ;
        RECT 0.060000 0.460000 0.130000 1.035000 ;
        RECT 0.425000 1.105000 0.560000 1.245000 ;
        RECT 0.995000 1.105000 1.130000 1.245000 ;
        RECT 1.755000 1.105000 1.890000 1.245000 ;
        RECT 0.060000 0.390000 0.750000 0.460000 ;
    END
    ANTENNADIFFAREA 0.3808 ;
    ANTENNAPARTIALMETALAREA 0.27335 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9321 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 0.085000 1.170000 0.155000 1.315000 ;
        RECT 0.835000 1.170000 0.905000 1.315000 ;
        RECT 1.405000 1.170000 1.475000 1.315000 ;
        RECT 1.975000 1.065000 2.045000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 1.185000 0.085000 1.320000 0.190000 ;
        RECT 1.565000 0.085000 1.700000 0.190000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.000000 0.390000 1.890000 0.460000 ;
      RECT 1.975000 0.325000 2.045000 0.425000 ;
      RECT 0.050000 0.255000 2.045000 0.325000 ;
      RECT 1.975000 0.150000 2.045000 0.255000 ;
  END
END OAI221_X2

MACRO OAI221_X4
  CLASS CORE ;
  FOREIGN OAI221_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.585000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.020125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0754 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.775000 0.525000 0.900000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.155000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.025375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.245000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.032375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0936 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.020125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0754 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.795000 0.185000 1.865000 0.700000 ;
        RECT 1.795000 0.700000 2.235000 0.840000 ;
        RECT 1.795000 0.840000 1.865000 1.250000 ;
        RECT 2.165000 0.840000 2.235000 1.250000 ;
        RECT 2.165000 0.185000 2.235000 0.700000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1911 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6318 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.470000 1.040000 0.540000 1.315000 ;
        RECT 1.190000 1.040000 1.260000 1.315000 ;
        RECT 1.595000 0.975000 1.665000 1.315000 ;
        RECT 1.975000 0.975000 2.045000 1.315000 ;
        RECT 2.355000 0.975000 2.425000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.820000 0.085000 0.955000 0.160000 ;
        RECT 1.190000 0.085000 1.260000 0.200000 ;
        RECT 1.595000 0.085000 1.665000 0.335000 ;
        RECT 1.975000 0.085000 2.045000 0.460000 ;
        RECT 2.355000 0.085000 2.425000 0.460000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.100000 0.220000 0.170000 0.285000 ;
      RECT 0.100000 0.150000 0.540000 0.220000 ;
      RECT 0.470000 0.220000 0.540000 0.285000 ;
      RECT 0.670000 0.255000 1.110000 0.325000 ;
      RECT 0.670000 0.150000 0.740000 0.255000 ;
      RECT 0.100000 0.845000 0.170000 1.120000 ;
      RECT 0.100000 0.775000 1.350000 0.845000 ;
      RECT 0.660000 0.845000 0.730000 1.120000 ;
      RECT 1.280000 0.460000 1.350000 0.775000 ;
      RECT 0.290000 0.390000 1.350000 0.460000 ;
      RECT 0.290000 0.285000 0.360000 0.390000 ;
      RECT 1.415000 0.660000 1.485000 1.250000 ;
      RECT 1.415000 0.525000 1.730000 0.660000 ;
      RECT 1.415000 0.185000 1.485000 0.525000 ;
  END
END OAI221_X4

MACRO OAI222_X1
  CLASS CORE ;
  FOREIGN OAI222_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.340000 0.525000 1.460000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.115000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.018375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.755000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.525000 0.945000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.350000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.028 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0871 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.200000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0819 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.520000 0.795000 1.430000 0.865000 ;
        RECT 0.520000 0.865000 0.590000 1.140000 ;
        RECT 1.360000 0.865000 1.430000 1.140000 ;
        RECT 1.180000 0.400000 1.270000 0.795000 ;
    END
    ANTENNADIFFAREA 0.3227 ;
    ANTENNAPARTIALMETALAREA 0.13775 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5005 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.520000 1.485000 ;
        RECT 0.050000 1.040000 0.120000 1.315000 ;
        RECT 0.980000 1.040000 1.050000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.520000 0.085000 ;
        RECT 0.050000 0.085000 0.120000 0.425000 ;
        RECT 0.395000 0.085000 0.530000 0.190000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.245000 0.325000 0.315000 0.425000 ;
      RECT 0.245000 0.255000 0.860000 0.325000 ;
      RECT 0.245000 0.150000 0.315000 0.255000 ;
      RECT 0.790000 0.150000 0.860000 0.255000 ;
      RECT 0.575000 0.390000 1.050000 0.460000 ;
      RECT 0.980000 0.335000 1.050000 0.390000 ;
      RECT 0.980000 0.265000 1.430000 0.335000 ;
      RECT 1.360000 0.335000 1.430000 0.425000 ;
      RECT 0.980000 0.150000 1.050000 0.265000 ;
      RECT 1.360000 0.150000 1.430000 0.265000 ;
  END
END OAI222_X1

MACRO OAI222_X2
  CLASS CORE ;
  FOREIGN OAI222_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.850000 0.525000 1.920000 0.725000 ;
        RECT 1.850000 0.725000 2.465000 0.795000 ;
        RECT 2.340000 0.525000 2.465000 0.725000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08205 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2821 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.150000 0.420000 2.220000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955000 0.525000 1.025000 0.770000 ;
        RECT 0.955000 0.770000 1.650000 0.840000 ;
        RECT 1.525000 0.525000 1.650000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.096425 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3263 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.200000 0.525000 1.290000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.320000 0.770000 ;
        RECT 0.195000 0.770000 0.830000 0.840000 ;
        RECT 0.760000 0.525000 0.830000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.092225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3107 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.530000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.090000 0.905000 2.600000 0.975000 ;
        RECT 0.090000 0.975000 0.160000 1.250000 ;
        RECT 0.840000 0.975000 0.910000 1.250000 ;
        RECT 1.605000 0.975000 1.675000 1.250000 ;
        RECT 2.530000 0.975000 2.600000 1.250000 ;
        RECT 2.530000 0.355000 2.600000 0.905000 ;
        RECT 1.925000 0.285000 2.600000 0.355000 ;
    END
    ANTENNADIFFAREA 0.52885 ;
    ANTENNAPARTIALMETALAREA 0.33845 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2753 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.660000 1.485000 ;
        RECT 0.460000 1.040000 0.530000 1.315000 ;
        RECT 1.220000 1.040000 1.290000 1.315000 ;
        RECT 2.140000 1.040000 2.210000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.660000 0.085000 ;
        RECT 0.270000 0.085000 0.340000 0.285000 ;
        RECT 0.650000 0.085000 0.720000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.090000 0.355000 0.910000 0.425000 ;
      RECT 0.840000 0.220000 0.910000 0.355000 ;
      RECT 0.090000 0.150000 0.160000 0.355000 ;
      RECT 0.465000 0.150000 0.535000 0.355000 ;
      RECT 0.840000 0.150000 1.705000 0.220000 ;
      RECT 1.005000 0.355000 1.840000 0.425000 ;
      RECT 1.770000 0.220000 1.840000 0.355000 ;
      RECT 1.770000 0.150000 2.625000 0.220000 ;
  END
END OAI222_X2

MACRO OAI222_X4
  CLASS CORE ;
  FOREIGN OAI222_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.560000 0.900000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.495000 0.560000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0287 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0897 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.560000 1.130000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.195000 0.560000 1.330000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.915000 0.150000 1.985000 0.560000 ;
        RECT 1.915000 0.560000 2.360000 0.700000 ;
        RECT 1.915000 0.700000 1.985000 1.250000 ;
        RECT 2.290000 0.700000 2.360000 1.250000 ;
        RECT 2.290000 0.150000 2.360000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1967 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6513 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.660000 1.485000 ;
        RECT 1.335000 1.040000 1.405000 1.315000 ;
        RECT 0.415000 1.030000 0.485000 1.315000 ;
        RECT 1.715000 0.975000 1.785000 1.315000 ;
        RECT 2.095000 0.975000 2.165000 1.315000 ;
        RECT 2.475000 0.975000 2.545000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.660000 0.085000 ;
        RECT 0.965000 0.085000 1.035000 0.220000 ;
        RECT 1.335000 0.085000 1.405000 0.220000 ;
        RECT 1.715000 0.085000 1.785000 0.335000 ;
        RECT 2.095000 0.085000 2.165000 0.425000 ;
        RECT 2.475000 0.085000 2.545000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.220000 0.115000 0.425000 ;
      RECT 0.045000 0.150000 0.900000 0.220000 ;
      RECT 0.580000 0.420000 1.250000 0.490000 ;
      RECT 0.045000 0.855000 0.115000 1.075000 ;
      RECT 0.045000 0.785000 1.465000 0.855000 ;
      RECT 0.880000 0.855000 0.950000 1.075000 ;
      RECT 1.395000 0.355000 1.465000 0.785000 ;
      RECT 0.200000 0.285000 1.465000 0.355000 ;
      RECT 1.535000 0.660000 1.605000 1.160000 ;
      RECT 1.535000 0.525000 1.850000 0.660000 ;
      RECT 1.535000 0.150000 1.605000 0.525000 ;
  END
END OAI222_X4

MACRO OAI22_X1
  CLASS CORE ;
  FOREIGN OAI22_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.390000 0.725000 0.460000 ;
        RECT 0.440000 0.460000 0.510000 1.050000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.06125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2457 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.055000 0.975000 0.125000 1.315000 ;
        RECT 0.810000 0.975000 0.880000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.210000 0.085000 0.345000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 0.315000 0.130000 0.460000 ;
      RECT 0.060000 0.245000 0.880000 0.315000 ;
      RECT 0.810000 0.315000 0.880000 0.460000 ;
      RECT 0.060000 0.185000 0.130000 0.245000 ;
      RECT 0.810000 0.185000 0.880000 0.245000 ;
  END
END OAI22_X1

MACRO OAI22_X2
  CLASS CORE ;
  FOREIGN OAI22_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.185000 0.525000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.525000 0.950000 0.765000 ;
        RECT 0.820000 0.765000 1.515000 0.835000 ;
        RECT 1.445000 0.525000 1.515000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09665 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3237 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.525000 0.525000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.765000 ;
        RECT 0.060000 0.765000 0.750000 0.835000 ;
        RECT 0.680000 0.525000 0.750000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0951 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3224 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.900000 1.650000 0.970000 ;
        RECT 0.425000 0.970000 0.495000 1.250000 ;
        RECT 1.185000 0.970000 1.255000 1.250000 ;
        RECT 1.580000 0.460000 1.650000 0.900000 ;
        RECT 0.960000 0.390000 1.650000 0.460000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.20405 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7761 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.040000 1.035000 0.110000 1.315000 ;
        RECT 0.795000 1.035000 0.865000 1.315000 ;
        RECT 1.555000 1.035000 1.625000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.355000 0.865000 0.425000 ;
      RECT 0.795000 0.220000 0.865000 0.355000 ;
      RECT 0.045000 0.150000 0.115000 0.355000 ;
      RECT 0.415000 0.150000 0.485000 0.355000 ;
      RECT 0.795000 0.150000 1.660000 0.220000 ;
  END
END OAI22_X2

MACRO DLL_X1
  CLASS CORE ;
  FOREIGN DLL_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.560000 0.430000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0252 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.580000 0.525000 1.705000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.390000 0.260000 1.460000 0.840000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0406 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.169 LAYER metal1 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.900000 1.485000 ;
        RECT 1.575000 1.040000 1.645000 1.315000 ;
        RECT 1.035000 0.950000 1.105000 1.315000 ;
        RECT 0.275000 0.915000 0.345000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.900000 0.085000 ;
        RECT 0.275000 0.085000 0.345000 0.415000 ;
        RECT 1.035000 0.085000 1.105000 0.420000 ;
        RECT 1.575000 0.085000 1.645000 0.235000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.095000 0.850000 0.165000 1.085000 ;
      RECT 0.095000 0.780000 0.600000 0.850000 ;
      RECT 0.530000 0.850000 0.600000 1.250000 ;
      RECT 0.095000 0.280000 0.165000 0.780000 ;
      RECT 0.530000 0.220000 0.600000 0.780000 ;
      RECT 0.530000 0.150000 0.845000 0.220000 ;
      RECT 0.665000 0.660000 0.735000 1.085000 ;
      RECT 0.665000 0.525000 1.165000 0.660000 ;
      RECT 0.665000 0.285000 0.735000 0.525000 ;
      RECT 1.230000 0.845000 1.300000 1.085000 ;
      RECT 0.900000 0.775000 1.300000 0.845000 ;
      RECT 1.230000 0.285000 1.300000 0.775000 ;
      RECT 1.235000 1.180000 1.510000 1.250000 ;
      RECT 1.440000 0.975000 1.510000 1.180000 ;
      RECT 1.440000 0.905000 1.840000 0.975000 ;
      RECT 1.770000 0.975000 1.840000 1.240000 ;
      RECT 1.770000 0.195000 1.840000 0.905000 ;
  END
END DLL_X1

MACRO DLL_X2
  CLASS CORE ;
  FOREIGN DLL_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.510000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0247 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.770000 0.525000 1.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END GN

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.580000 0.260000 1.650000 1.005000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.05215 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2119 LAYER metal1 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 1.385000 1.205000 1.455000 1.315000 ;
        RECT 1.760000 1.205000 1.830000 1.315000 ;
        RECT 0.225000 0.900000 0.295000 1.315000 ;
        RECT 0.985000 0.875000 1.055000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.370000 ;
        RECT 0.985000 0.085000 1.055000 0.460000 ;
        RECT 1.385000 0.085000 1.455000 0.395000 ;
        RECT 1.760000 0.085000 1.830000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.835000 0.115000 1.145000 ;
      RECT 0.045000 0.765000 0.550000 0.835000 ;
      RECT 0.045000 0.300000 0.115000 0.765000 ;
      RECT 0.480000 0.265000 0.550000 0.765000 ;
      RECT 0.480000 0.195000 0.820000 0.265000 ;
      RECT 0.615000 0.660000 0.685000 1.015000 ;
      RECT 0.615000 0.525000 1.125000 0.660000 ;
      RECT 0.615000 0.335000 0.685000 0.525000 ;
      RECT 1.190000 0.800000 1.260000 1.005000 ;
      RECT 0.850000 0.730000 1.260000 0.800000 ;
      RECT 1.190000 0.325000 1.260000 0.730000 ;
      RECT 1.185000 1.140000 1.320000 1.250000 ;
      RECT 1.185000 1.070000 2.025000 1.140000 ;
      RECT 1.955000 1.140000 2.025000 1.240000 ;
      RECT 1.955000 0.195000 2.025000 1.070000 ;
  END
END DLL_X2

MACRO FA_X1
  CLASS CORE ;
  FOREIGN FA_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.905000 0.825000 2.660000 0.895000 ;
        RECT 2.530000 0.700000 2.660000 0.825000 ;
    END
    ANTENNAGATEAREA 0.105 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1391 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.507 LAYER metal1 ;
    ANTENNAGATEAREA 0.105 LAYER metal2 ;
    ANTENNAGATEAREA 0.105 LAYER metal3 ;
    ANTENNAGATEAREA 0.105 LAYER metal4 ;
    ANTENNAGATEAREA 0.105 LAYER metal5 ;
    ANTENNAGATEAREA 0.105 LAYER metal6 ;
    ANTENNAGATEAREA 0.105 LAYER metal7 ;
    ANTENNAGATEAREA 0.105 LAYER metal8 ;
    ANTENNAGATEAREA 0.105 LAYER metal9 ;
    ANTENNAGATEAREA 0.105 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.410000 0.420000 2.470000 0.490000 ;
        RECT 2.340000 0.490000 2.470000 0.560000 ;
    END
    ANTENNAGATEAREA 0.105 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0833 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.312 LAYER metal1 ;
    ANTENNAGATEAREA 0.105 LAYER metal2 ;
    ANTENNAGATEAREA 0.105 LAYER metal3 ;
    ANTENNAGATEAREA 0.105 LAYER metal4 ;
    ANTENNAGATEAREA 0.105 LAYER metal5 ;
    ANTENNAGATEAREA 0.105 LAYER metal6 ;
    ANTENNAGATEAREA 0.105 LAYER metal7 ;
    ANTENNAGATEAREA 0.105 LAYER metal8 ;
    ANTENNAGATEAREA 0.105 LAYER metal9 ;
    ANTENNAGATEAREA 0.105 LAYER metal10 ;
  END B

  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.420000 0.700000 0.555000 ;
        RECT 0.630000 0.555000 2.275000 0.625000 ;
    END
    ANTENNAGATEAREA 0.07875 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1246 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.481 LAYER metal1 ;
    ANTENNAGATEAREA 0.07875 LAYER metal2 ;
    ANTENNAGATEAREA 0.07875 LAYER metal3 ;
    ANTENNAGATEAREA 0.07875 LAYER metal4 ;
    ANTENNAGATEAREA 0.07875 LAYER metal5 ;
    ANTENNAGATEAREA 0.07875 LAYER metal6 ;
    ANTENNAGATEAREA 0.07875 LAYER metal7 ;
    ANTENNAGATEAREA 0.07875 LAYER metal8 ;
    ANTENNAGATEAREA 0.07875 LAYER metal9 ;
    ANTENNAGATEAREA 0.07875 LAYER metal10 ;
  END CI

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.195000 0.135000 1.215000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0765 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2847 LAYER metal1 ;
  END CO

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.890000 0.195000 2.980000 1.215000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0918 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2886 LAYER metal1 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.040000 1.485000 ;
        RECT 2.695000 1.205000 2.765000 1.315000 ;
        RECT 1.015000 1.095000 1.085000 1.315000 ;
        RECT 1.705000 1.095000 1.840000 1.315000 ;
        RECT 1.360000 0.965000 1.430000 1.315000 ;
        RECT 0.250000 0.940000 0.320000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.040000 0.085000 ;
        RECT 0.250000 0.085000 0.320000 0.330000 ;
        RECT 1.025000 0.085000 1.095000 0.330000 ;
        RECT 1.360000 0.085000 1.430000 0.195000 ;
        RECT 1.705000 0.085000 1.840000 0.160000 ;
        RECT 2.665000 0.085000 2.800000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.835000 0.395000 1.275000 0.465000 ;
      RECT 0.835000 0.195000 0.905000 0.395000 ;
      RECT 1.205000 0.195000 1.275000 0.395000 ;
      RECT 0.800000 1.030000 0.935000 1.215000 ;
      RECT 0.800000 0.960000 1.275000 1.030000 ;
      RECT 1.205000 1.030000 1.275000 1.235000 ;
      RECT 1.555000 1.030000 1.625000 1.240000 ;
      RECT 1.555000 0.960000 2.000000 1.030000 ;
      RECT 1.930000 1.030000 2.000000 1.240000 ;
      RECT 1.520000 0.225000 2.030000 0.295000 ;
      RECT 0.630000 0.760000 0.700000 1.215000 ;
      RECT 0.495000 0.690000 2.115000 0.760000 ;
      RECT 0.495000 0.660000 0.565000 0.690000 ;
      RECT 0.205000 0.525000 0.565000 0.660000 ;
      RECT 0.495000 0.300000 0.565000 0.525000 ;
      RECT 0.495000 0.230000 0.735000 0.300000 ;
      RECT 2.130000 1.030000 2.200000 1.240000 ;
      RECT 2.130000 0.960000 2.820000 1.030000 ;
      RECT 2.750000 0.295000 2.820000 0.960000 ;
      RECT 2.100000 0.225000 2.820000 0.295000 ;
  END
END FA_X1

MACRO FILLCELL_X1
  CLASS CORE ;
  FOREIGN FILLCELL_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.190000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.190000 0.085000 ;
    END
  END VSS
END FILLCELL_X1

MACRO FILLCELL_X16
  CLASS CORE ;
  FOREIGN FILLCELL_X16 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.040000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.040000 0.085000 ;
    END
  END VSS
END FILLCELL_X16

MACRO FILLCELL_X2
  CLASS CORE ;
  FOREIGN FILLCELL_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.190000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.190000 0.085000 ;
    END
  END VSS
END FILLCELL_X2

MACRO FILLCELL_X32
  CLASS CORE ;
  FOREIGN FILLCELL_X32 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 6.08 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 6.080000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 6.080000 0.085000 ;
    END
  END VSS
END FILLCELL_X32

MACRO FILLCELL_X4
  CLASS CORE ;
  FOREIGN FILLCELL_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
    END
  END VSS
END FILLCELL_X4

MACRO FILLCELL_X8
  CLASS CORE ;
  FOREIGN FILLCELL_X8 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.520000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.520000 0.085000 ;
    END
  END VSS
END FILLCELL_X8

MACRO HA_X1
  CLASS CORE ;
  FOREIGN HA_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.355000 0.525000 0.425000 0.725000 ;
        RECT 0.355000 0.725000 0.740000 0.795000 ;
        RECT 0.670000 0.630000 0.740000 0.725000 ;
        RECT 0.670000 0.560000 1.080000 0.630000 ;
        RECT 1.010000 0.630000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.10475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0812 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3198 LAYER metal1 ;
    ANTENNAGATEAREA 0.10475 LAYER metal2 ;
    ANTENNAGATEAREA 0.10475 LAYER metal3 ;
    ANTENNAGATEAREA 0.10475 LAYER metal4 ;
    ANTENNAGATEAREA 0.10475 LAYER metal5 ;
    ANTENNAGATEAREA 0.10475 LAYER metal6 ;
    ANTENNAGATEAREA 0.10475 LAYER metal7 ;
    ANTENNAGATEAREA 0.10475 LAYER metal8 ;
    ANTENNAGATEAREA 0.10475 LAYER metal9 ;
    ANTENNAGATEAREA 0.10475 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.265000 0.860000 ;
        RECT 0.195000 0.860000 0.890000 0.930000 ;
        RECT 0.805000 0.700000 0.890000 0.860000 ;
    END
    ANTENNAGATEAREA 0.10475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0857 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3276 LAYER metal1 ;
    ANTENNAGATEAREA 0.10475 LAYER metal2 ;
    ANTENNAGATEAREA 0.10475 LAYER metal3 ;
    ANTENNAGATEAREA 0.10475 LAYER metal4 ;
    ANTENNAGATEAREA 0.10475 LAYER metal5 ;
    ANTENNAGATEAREA 0.10475 LAYER metal6 ;
    ANTENNAGATEAREA 0.10475 LAYER metal7 ;
    ANTENNAGATEAREA 0.10475 LAYER metal8 ;
    ANTENNAGATEAREA 0.10475 LAYER metal9 ;
    ANTENNAGATEAREA 0.10475 LAYER metal10 ;
  END B

  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.770000 0.150000 1.850000 1.250000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.088 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3068 LAYER metal1 ;
  END CO

  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.290000 0.525000 0.360000 ;
        RECT 0.060000 0.360000 0.130000 0.995000 ;
        RECT 0.455000 0.150000 0.525000 0.290000 ;
        RECT 0.060000 0.995000 0.370000 1.065000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.1085 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4212 LAYER metal1 ;
  END S

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.900000 1.485000 ;
        RECT 0.645000 1.080000 0.715000 1.315000 ;
        RECT 1.590000 1.080000 1.660000 1.315000 ;
        RECT 1.220000 0.940000 1.290000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.900000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.225000 ;
        RECT 0.645000 0.085000 0.715000 0.285000 ;
        RECT 1.030000 0.085000 1.100000 0.285000 ;
        RECT 1.590000 0.085000 1.660000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.050000 1.130000 0.560000 1.200000 ;
      RECT 1.035000 0.835000 1.105000 1.115000 ;
      RECT 1.035000 0.765000 1.250000 0.835000 ;
      RECT 1.180000 0.495000 1.250000 0.765000 ;
      RECT 0.535000 0.425000 1.250000 0.495000 ;
      RECT 0.535000 0.495000 0.605000 0.660000 ;
      RECT 0.840000 0.150000 0.910000 0.425000 ;
      RECT 1.400000 0.660000 1.470000 1.115000 ;
      RECT 1.400000 0.525000 1.705000 0.660000 ;
      RECT 1.400000 0.285000 1.470000 0.525000 ;
      RECT 1.220000 0.150000 1.470000 0.285000 ;
  END
END HA_X1

MACRO INV_X1
  CLASS CORE ;
  FOREIGN INV_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.165000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.018375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.230000 0.150000 0.325000 1.250000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3107 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.380000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.380000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
    END
  END VSS
END INV_X1

MACRO INV_X16
  CLASS CORE ;
  FOREIGN INV_X16 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.095000 0.525000 0.165000 1.050000 ;
        RECT 0.095000 1.050000 3.095000 1.120000 ;
        RECT 1.200000 0.525000 1.270000 1.050000 ;
        RECT 2.000000 0.525000 2.070000 1.050000 ;
        RECT 3.025000 0.525000 3.095000 1.050000 ;
    END
    ANTENNAGATEAREA 0.836 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.357 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3442 LAYER metal1 ;
    ANTENNAGATEAREA 0.836 LAYER metal2 ;
    ANTENNAGATEAREA 0.836 LAYER metal3 ;
    ANTENNAGATEAREA 0.836 LAYER metal4 ;
    ANTENNAGATEAREA 0.836 LAYER metal5 ;
    ANTENNAGATEAREA 0.836 LAYER metal6 ;
    ANTENNAGATEAREA 0.836 LAYER metal7 ;
    ANTENNAGATEAREA 0.836 LAYER metal8 ;
    ANTENNAGATEAREA 0.836 LAYER metal9 ;
    ANTENNAGATEAREA 0.836 LAYER metal10 ;
  END A

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.180000 0.305000 0.280000 ;
        RECT 0.235000 0.280000 2.955000 0.420000 ;
        RECT 0.235000 0.420000 0.305000 0.985000 ;
        RECT 0.605000 0.420000 0.675000 0.985000 ;
        RECT 0.985000 0.420000 1.055000 0.985000 ;
        RECT 1.365000 0.420000 1.435000 0.985000 ;
        RECT 1.745000 0.420000 1.815000 0.985000 ;
        RECT 2.135000 0.420000 2.205000 0.985000 ;
        RECT 2.505000 0.420000 2.575000 0.985000 ;
        RECT 2.885000 0.420000 2.955000 0.985000 ;
        RECT 0.605000 0.160000 0.675000 0.280000 ;
        RECT 0.985000 0.150000 1.055000 0.280000 ;
        RECT 1.365000 0.150000 1.435000 0.280000 ;
        RECT 1.745000 0.150000 1.815000 0.280000 ;
        RECT 2.125000 0.150000 2.195000 0.280000 ;
        RECT 2.505000 0.150000 2.575000 0.280000 ;
        RECT 2.885000 0.150000 2.955000 0.280000 ;
    END
    ANTENNADIFFAREA 1.1704 ;
    ANTENNAPARTIALMETALAREA 0.7672 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1788 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.230000 1.485000 ;
        RECT 0.040000 1.205000 0.110000 1.315000 ;
        RECT 0.415000 1.205000 0.485000 1.315000 ;
        RECT 0.795000 1.205000 0.865000 1.315000 ;
        RECT 1.175000 1.205000 1.245000 1.315000 ;
        RECT 1.555000 1.205000 1.625000 1.315000 ;
        RECT 1.935000 1.205000 2.005000 1.315000 ;
        RECT 2.315000 1.205000 2.385000 1.315000 ;
        RECT 2.695000 1.205000 2.765000 1.315000 ;
        RECT 3.075000 1.205000 3.145000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.230000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.365000 ;
        RECT 0.415000 0.085000 0.485000 0.210000 ;
        RECT 0.795000 0.085000 0.865000 0.210000 ;
        RECT 1.175000 0.085000 1.245000 0.210000 ;
        RECT 1.555000 0.085000 1.625000 0.210000 ;
        RECT 1.935000 0.085000 2.005000 0.210000 ;
        RECT 2.315000 0.085000 2.385000 0.210000 ;
        RECT 2.695000 0.085000 2.765000 0.210000 ;
        RECT 3.075000 0.085000 3.145000 0.365000 ;
    END
  END VSS
END INV_X16

MACRO INV_X2
  CLASS CORE ;
  FOREIGN INV_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.150000 0.320000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.077 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3042 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.570000 1.485000 ;
        RECT 0.055000 0.975000 0.125000 1.315000 ;
        RECT 0.430000 0.975000 0.500000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.570000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.425000 ;
        RECT 0.430000 0.085000 0.500000 0.425000 ;
    END
  END VSS
END INV_X2

MACRO INV_X32
  CLASS CORE ;
  FOREIGN INV_X32 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 6.27 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.115000 0.525000 0.185000 0.930000 ;
        RECT 0.115000 0.930000 5.850000 1.000000 ;
        RECT 1.200000 0.525000 1.270000 0.930000 ;
        RECT 2.340000 0.525000 2.410000 0.930000 ;
        RECT 3.480000 0.525000 3.550000 0.930000 ;
        RECT 4.620000 0.525000 4.690000 0.930000 ;
        RECT 5.780000 0.525000 5.850000 0.930000 ;
    END
    ANTENNAGATEAREA 1.672 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.57155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1411 LAYER metal1 ;
    ANTENNAGATEAREA 1.672 LAYER metal2 ;
    ANTENNAGATEAREA 1.672 LAYER metal3 ;
    ANTENNAGATEAREA 1.672 LAYER metal4 ;
    ANTENNAGATEAREA 1.672 LAYER metal5 ;
    ANTENNAGATEAREA 1.672 LAYER metal6 ;
    ANTENNAGATEAREA 1.672 LAYER metal7 ;
    ANTENNAGATEAREA 1.672 LAYER metal8 ;
    ANTENNAGATEAREA 1.672 LAYER metal9 ;
    ANTENNAGATEAREA 1.672 LAYER metal10 ;
  END A

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.160000 0.320000 0.280000 ;
        RECT 0.250000 0.280000 6.015000 0.420000 ;
        RECT 0.250000 0.420000 0.320000 0.865000 ;
        RECT 0.620000 0.420000 0.690000 0.865000 ;
        RECT 1.000000 0.420000 1.070000 0.865000 ;
        RECT 1.390000 0.420000 1.460000 0.865000 ;
        RECT 1.760000 0.420000 1.830000 0.865000 ;
        RECT 2.140000 0.420000 2.210000 0.865000 ;
        RECT 2.525000 0.420000 2.595000 0.865000 ;
        RECT 2.900000 0.420000 2.970000 0.865000 ;
        RECT 3.280000 0.420000 3.350000 0.865000 ;
        RECT 3.665000 0.420000 3.735000 0.865000 ;
        RECT 4.040000 0.420000 4.110000 0.865000 ;
        RECT 4.420000 0.420000 4.490000 0.865000 ;
        RECT 4.810000 0.420000 4.880000 0.865000 ;
        RECT 5.180000 0.420000 5.250000 0.865000 ;
        RECT 5.560000 0.420000 5.630000 0.865000 ;
        RECT 5.945000 0.420000 6.015000 1.005000 ;
        RECT 0.620000 0.160000 0.690000 0.280000 ;
        RECT 1.000000 0.160000 1.070000 0.280000 ;
        RECT 1.390000 0.160000 1.460000 0.280000 ;
        RECT 1.760000 0.160000 1.830000 0.280000 ;
        RECT 2.140000 0.160000 2.210000 0.280000 ;
        RECT 2.525000 0.160000 2.595000 0.280000 ;
        RECT 2.900000 0.160000 2.970000 0.280000 ;
        RECT 3.280000 0.160000 3.350000 0.280000 ;
        RECT 3.665000 0.160000 3.735000 0.280000 ;
        RECT 4.040000 0.160000 4.110000 0.280000 ;
        RECT 4.420000 0.160000 4.490000 0.280000 ;
        RECT 4.800000 0.160000 4.870000 0.280000 ;
        RECT 5.180000 0.160000 5.250000 0.280000 ;
        RECT 5.560000 0.160000 5.630000 0.280000 ;
        RECT 5.945000 0.160000 6.015000 0.280000 ;
    END
    ANTENNADIFFAREA 2.3408 ;
    ANTENNAPARTIALMETALAREA 1.4497 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.9221 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 6.270000 1.485000 ;
        RECT 0.055000 1.065000 0.125000 1.315000 ;
        RECT 0.430000 1.065000 0.500000 1.315000 ;
        RECT 0.810000 1.065000 0.880000 1.315000 ;
        RECT 1.190000 1.065000 1.260000 1.315000 ;
        RECT 1.570000 1.065000 1.640000 1.315000 ;
        RECT 1.950000 1.065000 2.020000 1.315000 ;
        RECT 2.330000 1.065000 2.400000 1.315000 ;
        RECT 2.710000 1.065000 2.780000 1.315000 ;
        RECT 3.090000 1.065000 3.160000 1.315000 ;
        RECT 3.470000 1.065000 3.540000 1.315000 ;
        RECT 3.850000 1.065000 3.920000 1.315000 ;
        RECT 4.230000 1.065000 4.300000 1.315000 ;
        RECT 4.610000 1.065000 4.680000 1.315000 ;
        RECT 4.990000 1.065000 5.060000 1.315000 ;
        RECT 5.370000 1.065000 5.440000 1.315000 ;
        RECT 5.750000 1.065000 5.820000 1.315000 ;
        RECT 6.130000 1.065000 6.200000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 6.270000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.335000 ;
        RECT 0.430000 0.085000 0.500000 0.195000 ;
        RECT 0.810000 0.085000 0.880000 0.195000 ;
        RECT 1.190000 0.085000 1.260000 0.195000 ;
        RECT 1.570000 0.085000 1.640000 0.195000 ;
        RECT 1.950000 0.085000 2.020000 0.195000 ;
        RECT 2.330000 0.085000 2.400000 0.195000 ;
        RECT 2.710000 0.085000 2.780000 0.195000 ;
        RECT 3.090000 0.085000 3.160000 0.195000 ;
        RECT 3.470000 0.085000 3.540000 0.195000 ;
        RECT 3.850000 0.085000 3.920000 0.195000 ;
        RECT 4.230000 0.085000 4.300000 0.195000 ;
        RECT 4.610000 0.085000 4.680000 0.195000 ;
        RECT 4.990000 0.085000 5.060000 0.195000 ;
        RECT 5.370000 0.085000 5.440000 0.195000 ;
        RECT 5.750000 0.085000 5.820000 0.195000 ;
        RECT 6.130000 0.085000 6.200000 0.335000 ;
    END
  END VSS
END INV_X32

MACRO INV_X4
  CLASS CORE ;
  FOREIGN INV_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.170000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.150000 0.305000 0.560000 ;
        RECT 0.235000 0.560000 0.685000 0.700000 ;
        RECT 0.235000 0.700000 0.305000 1.040000 ;
        RECT 0.615000 0.700000 0.685000 1.040000 ;
        RECT 0.610000 0.150000 0.685000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.17005 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5434 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.040000 0.980000 0.110000 1.315000 ;
        RECT 0.415000 0.980000 0.485000 1.315000 ;
        RECT 0.795000 0.980000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.425000 ;
        RECT 0.795000 0.085000 0.865000 0.425000 ;
    END
  END VSS
END INV_X4

MACRO INV_X8
  CLASS CORE ;
  FOREIGN INV_X8 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.170000 0.700000 ;
    END
    ANTENNAGATEAREA 0.418 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.418 LAYER metal2 ;
    ANTENNAGATEAREA 0.418 LAYER metal3 ;
    ANTENNAGATEAREA 0.418 LAYER metal4 ;
    ANTENNAGATEAREA 0.418 LAYER metal5 ;
    ANTENNAGATEAREA 0.418 LAYER metal6 ;
    ANTENNAGATEAREA 0.418 LAYER metal7 ;
    ANTENNAGATEAREA 0.418 LAYER metal8 ;
    ANTENNAGATEAREA 0.418 LAYER metal9 ;
    ANTENNAGATEAREA 0.418 LAYER metal10 ;
  END A

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.150000 0.305000 0.560000 ;
        RECT 0.235000 0.560000 1.445000 0.700000 ;
        RECT 0.235000 0.700000 0.305000 1.040000 ;
        RECT 0.605000 0.700000 0.675000 1.040000 ;
        RECT 0.985000 0.700000 1.055000 1.040000 ;
        RECT 1.375000 0.700000 1.445000 1.040000 ;
        RECT 0.605000 0.150000 0.675000 0.560000 ;
        RECT 0.985000 0.150000 1.055000 0.560000 ;
        RECT 1.375000 0.150000 1.445000 0.560000 ;
    END
    ANTENNADIFFAREA 0.5852 ;
    ANTENNAPARTIALMETALAREA 0.3794 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.131 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.040000 0.970000 0.110000 1.315000 ;
        RECT 0.415000 0.970000 0.485000 1.315000 ;
        RECT 0.795000 0.970000 0.865000 1.315000 ;
        RECT 1.175000 0.970000 1.245000 1.315000 ;
        RECT 1.555000 0.970000 1.625000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.360000 ;
        RECT 0.415000 0.085000 0.485000 0.360000 ;
        RECT 0.795000 0.085000 0.865000 0.360000 ;
        RECT 1.175000 0.085000 1.245000 0.360000 ;
        RECT 1.555000 0.085000 1.625000 0.360000 ;
    END
  END VSS
END INV_X8

MACRO LOGIC0_X1
  CLASS CORE ;
  FOREIGN LOGIC0_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.150000 0.130000 0.840000 ;
    END
    ANTENNADIFFAREA 0.00945 ;
    ANTENNAPARTIALMETALAREA 0.0483 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1976 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.380000 1.485000 ;
        RECT 0.245000 1.115000 0.315000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.380000 0.085000 ;
        RECT 0.240000 0.085000 0.310000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 0.975000 0.180000 1.250000 ;
  END
END LOGIC0_X1

MACRO LOGIC1_X1
  CLASS CORE ;
  FOREIGN LOGIC1_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.38 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.560000 0.130000 1.250000 ;
    END
    ANTENNADIFFAREA 0.014175 ;
    ANTENNAPARTIALMETALAREA 0.0483 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1976 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.380000 1.485000 ;
        RECT 0.240000 1.115000 0.310000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.380000 0.085000 ;
        RECT 0.245000 0.085000 0.315000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 0.150000 0.180000 0.425000 ;
  END
END LOGIC1_X1

MACRO MUX2_X1
  CLASS CORE ;
  FOREIGN MUX2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.525000 0.950000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END B

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.765000 ;
        RECT 0.060000 0.765000 0.595000 0.835000 ;
        RECT 0.525000 0.535000 0.595000 0.765000 ;
    END
    ANTENNAGATEAREA 0.0525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08355 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2795 LAYER metal1 ;
    ANTENNAGATEAREA 0.0525 LAYER metal2 ;
    ANTENNAGATEAREA 0.0525 LAYER metal3 ;
    ANTENNAGATEAREA 0.0525 LAYER metal4 ;
    ANTENNAGATEAREA 0.0525 LAYER metal5 ;
    ANTENNAGATEAREA 0.0525 LAYER metal6 ;
    ANTENNAGATEAREA 0.0525 LAYER metal7 ;
    ANTENNAGATEAREA 0.0525 LAYER metal8 ;
    ANTENNAGATEAREA 0.0525 LAYER metal9 ;
    ANTENNAGATEAREA 0.0525 LAYER metal10 ;
  END S

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.180000 0.190000 1.270000 1.230000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0936 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2938 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.225000 1.035000 0.295000 1.315000 ;
        RECT 0.985000 0.975000 1.055000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.240000 ;
        RECT 0.985000 0.085000 1.055000 0.240000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.970000 0.115000 1.250000 ;
      RECT 0.045000 0.900000 0.755000 0.970000 ;
      RECT 0.685000 0.460000 0.755000 0.900000 ;
      RECT 0.045000 0.390000 0.755000 0.460000 ;
      RECT 0.045000 0.190000 0.115000 0.390000 ;
      RECT 0.580000 1.070000 0.920000 1.140000 ;
      RECT 0.850000 0.910000 0.920000 1.070000 ;
      RECT 0.850000 0.840000 1.115000 0.910000 ;
      RECT 1.045000 0.460000 1.115000 0.840000 ;
      RECT 0.830000 0.390000 1.115000 0.460000 ;
      RECT 0.830000 0.290000 0.900000 0.390000 ;
      RECT 0.580000 0.220000 0.900000 0.290000 ;
  END
END MUX2_X1

MACRO MUX2_X2
  CLASS CORE ;
  FOREIGN MUX2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.225000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.028875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0884 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B

  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.770000 0.525000 0.995000 0.700000 ;
        RECT 0.925000 0.700000 0.995000 0.850000 ;
        RECT 0.925000 0.850000 1.535000 0.920000 ;
        RECT 1.465000 0.525000 1.535000 0.850000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.115325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3861 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END S

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.200000 0.150000 1.290000 0.785000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.05715 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1885 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.240000 1.240000 0.375000 1.315000 ;
        RECT 1.035000 1.205000 1.105000 1.315000 ;
        RECT 1.405000 1.205000 1.475000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.460000 0.085000 0.530000 0.285000 ;
        RECT 1.030000 0.085000 1.100000 0.285000 ;
        RECT 1.405000 0.085000 1.475000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.460000 1.175000 0.955000 1.245000 ;
      RECT 0.460000 1.135000 0.530000 1.175000 ;
      RECT 0.090000 1.065000 0.530000 1.135000 ;
      RECT 0.090000 0.860000 0.160000 1.065000 ;
      RECT 0.655000 0.970000 0.725000 1.075000 ;
      RECT 0.290000 0.900000 0.725000 0.970000 ;
      RECT 0.290000 0.455000 0.360000 0.900000 ;
      RECT 0.090000 0.385000 1.135000 0.455000 ;
      RECT 1.065000 0.455000 1.135000 0.660000 ;
      RECT 0.090000 0.150000 0.160000 0.385000 ;
      RECT 0.845000 0.150000 0.915000 0.385000 ;
      RECT 1.600000 1.055000 1.670000 1.250000 ;
      RECT 0.790000 0.985000 1.670000 1.055000 ;
      RECT 0.790000 0.835000 0.860000 0.985000 ;
      RECT 1.600000 0.150000 1.670000 0.985000 ;
      RECT 0.425000 0.765000 0.860000 0.835000 ;
      RECT 0.425000 0.525000 0.495000 0.765000 ;
  END
END MUX2_X2

MACRO NAND2_X1
  CLASS CORE ;
  FOREIGN NAND2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.355000 0.500000 0.425000 ;
        RECT 0.250000 0.425000 0.320000 1.250000 ;
        RECT 0.430000 0.150000 0.500000 0.355000 ;
    END
    ANTENNADIFFAREA 0.131775 ;
    ANTENNAPARTIALMETALAREA 0.0896 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.351 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.570000 1.485000 ;
        RECT 0.055000 0.975000 0.125000 1.315000 ;
        RECT 0.430000 0.975000 0.500000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.570000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.425000 ;
    END
  END VSS
END NAND2_X1

MACRO NAND2_X2
  CLASS CORE ;
  FOREIGN NAND2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0637 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.175000 0.525000 0.320000 0.660000 ;
        RECT 0.250000 0.660000 0.320000 0.770000 ;
        RECT 0.250000 0.770000 0.810000 0.840000 ;
        RECT 0.740000 0.525000 0.810000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.083625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3107 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.040000 0.460000 0.110000 0.905000 ;
        RECT 0.040000 0.905000 0.700000 0.975000 ;
        RECT 0.040000 0.390000 0.510000 0.460000 ;
        RECT 0.250000 0.975000 0.320000 1.250000 ;
        RECT 0.630000 0.975000 0.700000 1.250000 ;
        RECT 0.440000 0.150000 0.510000 0.390000 ;
    END
    ANTENNADIFFAREA 0.2345 ;
    ANTENNAPARTIALMETALAREA 0.16555 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6331 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.065000 1.040000 0.135000 1.315000 ;
        RECT 0.440000 1.040000 0.510000 1.315000 ;
        RECT 0.820000 1.040000 0.890000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.065000 0.085000 0.135000 0.285000 ;
        RECT 0.820000 0.085000 0.890000 0.425000 ;
    END
  END VSS
END NAND2_X2

MACRO NAND2_X4
  CLASS CORE ;
  FOREIGN NAND2_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.140000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.380000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.275000 0.785000 1.475000 0.855000 ;
        RECT 0.275000 0.855000 0.345000 1.070000 ;
        RECT 0.645000 0.855000 0.715000 1.070000 ;
        RECT 1.025000 0.855000 1.095000 1.070000 ;
        RECT 1.405000 0.855000 1.475000 1.070000 ;
        RECT 1.390000 0.420000 1.475000 0.785000 ;
        RECT 1.000000 0.350000 1.475000 0.420000 ;
    END
    ANTENNADIFFAREA 0.469 ;
    ANTENNAPARTIALMETALAREA 0.208475 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7683 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.080000 1.040000 0.150000 1.315000 ;
        RECT 0.455000 1.040000 0.525000 1.315000 ;
        RECT 0.835000 1.040000 0.905000 1.315000 ;
        RECT 1.215000 1.040000 1.285000 1.315000 ;
        RECT 1.595000 1.040000 1.665000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.265000 0.085000 0.335000 0.285000 ;
        RECT 0.645000 0.085000 0.715000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085000 0.355000 0.905000 0.425000 ;
      RECT 0.835000 0.220000 0.905000 0.355000 ;
      RECT 0.085000 0.150000 0.155000 0.355000 ;
      RECT 0.455000 0.150000 0.525000 0.355000 ;
      RECT 0.835000 0.150000 1.665000 0.220000 ;
      RECT 1.595000 0.220000 1.665000 0.425000 ;
  END
END NAND2_X4

MACRO NAND3_X1
  CLASS CORE ;
  FOREIGN NAND3_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.540000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.235000 0.800000 0.675000 0.870000 ;
        RECT 0.235000 0.870000 0.320000 1.250000 ;
        RECT 0.605000 0.870000 0.675000 1.250000 ;
        RECT 0.605000 0.150000 0.675000 0.800000 ;
    END
    ANTENNADIFFAREA 0.197925 ;
    ANTENNAPARTIALMETALAREA 0.1352 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4992 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
    END
  END VSS
END NAND3_X1

MACRO NAND3_X2
  CLASS CORE ;
  FOREIGN NAND3_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.595000 0.560000 0.730000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.380000 0.420000 1.080000 0.490000 ;
        RECT 0.380000 0.490000 0.450000 0.660000 ;
        RECT 0.950000 0.490000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0882 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.299 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.525000 0.265000 0.700000 ;
        RECT 0.195000 0.700000 0.320000 0.770000 ;
        RECT 0.195000 0.770000 1.215000 0.840000 ;
        RECT 1.145000 0.525000 1.215000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.10955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4108 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.335000 0.130000 0.905000 ;
        RECT 0.060000 0.905000 1.095000 0.975000 ;
        RECT 0.060000 0.265000 0.750000 0.335000 ;
        RECT 0.265000 0.975000 0.335000 1.250000 ;
        RECT 0.645000 0.975000 0.715000 1.250000 ;
        RECT 1.025000 0.975000 1.095000 1.250000 ;
    END
    ANTENNADIFFAREA 0.3227 ;
    ANTENNAPARTIALMETALAREA 0.2184 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8294 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.080000 1.040000 0.150000 1.315000 ;
        RECT 0.455000 1.040000 0.525000 1.315000 ;
        RECT 0.835000 1.040000 0.905000 1.315000 ;
        RECT 1.215000 1.040000 1.285000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.195000 ;
        RECT 1.215000 0.085000 1.285000 0.335000 ;
    END
  END VSS
END NAND3_X2

MACRO NAND3_X4
  CLASS CORE ;
  FOREIGN NAND3_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.625000 0.555000 0.890000 0.625000 ;
        RECT 0.820000 0.360000 0.890000 0.555000 ;
        RECT 0.820000 0.290000 1.730000 0.360000 ;
        RECT 1.660000 0.360000 1.730000 0.555000 ;
        RECT 1.660000 0.555000 1.890000 0.625000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.12565 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4849 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.380000 0.525000 0.450000 0.690000 ;
        RECT 0.380000 0.690000 1.080000 0.760000 ;
        RECT 0.955000 0.495000 1.080000 0.690000 ;
        RECT 0.955000 0.425000 1.595000 0.495000 ;
        RECT 1.525000 0.495000 1.595000 0.690000 ;
        RECT 1.525000 0.690000 2.130000 0.760000 ;
        RECT 2.060000 0.525000 2.130000 0.690000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.197275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6968 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.190000 0.525000 0.260000 0.825000 ;
        RECT 0.190000 0.825000 2.300000 0.895000 ;
        RECT 1.190000 0.560000 1.325000 0.825000 ;
        RECT 2.230000 0.525000 2.300000 0.825000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.225475 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7917 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.055000 0.425000 0.125000 0.980000 ;
        RECT 0.055000 0.980000 2.435000 1.050000 ;
        RECT 0.055000 0.355000 0.715000 0.425000 ;
        RECT 0.265000 1.050000 2.235000 1.120000 ;
        RECT 2.365000 0.425000 2.435000 0.980000 ;
        RECT 0.645000 0.150000 0.715000 0.355000 ;
        RECT 0.265000 1.120000 0.335000 1.220000 ;
        RECT 0.645000 1.120000 0.715000 1.220000 ;
        RECT 1.025000 1.120000 1.095000 1.220000 ;
        RECT 1.405000 1.120000 1.475000 1.220000 ;
        RECT 1.785000 1.120000 1.855000 1.220000 ;
        RECT 2.165000 1.120000 2.235000 1.220000 ;
        RECT 1.795000 0.355000 2.435000 0.425000 ;
        RECT 1.795000 0.150000 1.865000 0.355000 ;
    END
    ANTENNADIFFAREA 0.6454 ;
    ANTENNAPARTIALMETALAREA 0.5439 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5444 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 1.185000 1.205000 1.320000 1.315000 ;
        RECT 1.565000 1.205000 1.700000 1.315000 ;
        RECT 1.945000 1.205000 2.080000 1.315000 ;
        RECT 0.425000 1.195000 0.560000 1.315000 ;
        RECT 0.805000 1.195000 0.940000 1.315000 ;
        RECT 2.355000 1.170000 2.425000 1.315000 ;
        RECT 0.080000 1.160000 0.150000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.195000 ;
        RECT 1.215000 0.085000 1.285000 0.195000 ;
        RECT 2.355000 0.085000 2.425000 0.195000 ;
    END
  END VSS
END NAND3_X4

MACRO BUF_X16
  CLASS CORE ;
  FOREIGN BUF_X16 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.75 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.715000 ;
    END
    ANTENNAGATEAREA 0.418 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0819 LAYER metal1 ;
    ANTENNAGATEAREA 0.418 LAYER metal2 ;
    ANTENNAGATEAREA 0.418 LAYER metal3 ;
    ANTENNAGATEAREA 0.418 LAYER metal4 ;
    ANTENNAGATEAREA 0.418 LAYER metal5 ;
    ANTENNAGATEAREA 0.418 LAYER metal6 ;
    ANTENNAGATEAREA 0.418 LAYER metal7 ;
    ANTENNAGATEAREA 0.418 LAYER metal8 ;
    ANTENNAGATEAREA 0.418 LAYER metal9 ;
    ANTENNAGATEAREA 0.418 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.770000 0.150000 1.840000 0.280000 ;
        RECT 1.770000 0.280000 4.490000 0.420000 ;
        RECT 1.770000 0.420000 1.840000 0.925000 ;
        RECT 2.140000 0.420000 2.210000 0.925000 ;
        RECT 2.520000 0.420000 2.590000 0.925000 ;
        RECT 2.900000 0.420000 2.970000 0.925000 ;
        RECT 3.280000 0.420000 3.350000 0.925000 ;
        RECT 3.660000 0.420000 3.730000 0.925000 ;
        RECT 4.050000 0.420000 4.120000 0.925000 ;
        RECT 4.420000 0.420000 4.490000 0.925000 ;
        RECT 2.140000 0.150000 2.210000 0.280000 ;
        RECT 2.520000 0.150000 2.590000 0.280000 ;
        RECT 2.900000 0.150000 2.970000 0.280000 ;
        RECT 3.280000 0.150000 3.350000 0.280000 ;
        RECT 3.660000 0.150000 3.730000 0.280000 ;
        RECT 4.040000 0.150000 4.110000 0.280000 ;
        RECT 4.420000 0.150000 4.490000 0.280000 ;
    END
    ANTENNADIFFAREA 1.1704 ;
    ANTENNAPARTIALMETALAREA 0.7364 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0644 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.750000 1.485000 ;
        RECT 1.570000 1.205000 1.640000 1.315000 ;
        RECT 1.950000 1.205000 2.020000 1.315000 ;
        RECT 2.330000 1.205000 2.400000 1.315000 ;
        RECT 2.710000 1.205000 2.780000 1.315000 ;
        RECT 3.090000 1.205000 3.160000 1.315000 ;
        RECT 3.470000 1.205000 3.540000 1.315000 ;
        RECT 3.850000 1.205000 3.920000 1.315000 ;
        RECT 4.230000 1.205000 4.300000 1.315000 ;
        RECT 4.610000 1.205000 4.680000 1.315000 ;
        RECT 0.055000 0.975000 0.125000 1.315000 ;
        RECT 0.430000 0.975000 0.500000 1.315000 ;
        RECT 0.810000 0.975000 0.880000 1.315000 ;
        RECT 1.190000 0.975000 1.260000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.750000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.340000 ;
        RECT 0.430000 0.085000 0.500000 0.340000 ;
        RECT 0.810000 0.085000 0.880000 0.340000 ;
        RECT 1.190000 0.085000 1.260000 0.340000 ;
        RECT 1.570000 0.085000 1.640000 0.340000 ;
        RECT 1.950000 0.085000 2.020000 0.200000 ;
        RECT 2.330000 0.085000 2.400000 0.200000 ;
        RECT 2.710000 0.085000 2.780000 0.200000 ;
        RECT 3.090000 0.085000 3.160000 0.200000 ;
        RECT 3.470000 0.085000 3.540000 0.200000 ;
        RECT 3.850000 0.085000 3.920000 0.200000 ;
        RECT 4.230000 0.085000 4.300000 0.200000 ;
        RECT 4.610000 0.085000 4.680000 0.200000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.250000 0.660000 0.320000 1.250000 ;
      RECT 0.250000 0.525000 1.705000 0.660000 ;
      RECT 0.620000 0.660000 0.690000 1.250000 ;
      RECT 1.000000 0.660000 1.070000 1.250000 ;
      RECT 1.380000 0.660000 1.450000 1.250000 ;
      RECT 1.635000 0.660000 1.705000 1.050000 ;
      RECT 0.250000 0.150000 0.320000 0.525000 ;
      RECT 0.620000 0.150000 0.690000 0.525000 ;
      RECT 1.000000 0.150000 1.070000 0.525000 ;
      RECT 1.380000 0.150000 1.450000 0.525000 ;
      RECT 1.635000 1.050000 4.630000 1.120000 ;
      RECT 2.690000 0.525000 2.760000 1.050000 ;
      RECT 3.450000 0.525000 3.520000 1.050000 ;
      RECT 4.560000 0.525000 4.630000 1.050000 ;
  END
END BUF_X16

MACRO BUF_X2
  CLASS CORE ;
  FOREIGN BUF_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.230000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0897 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.465000 0.150000 0.535000 0.560000 ;
        RECT 0.465000 0.560000 0.700000 0.700000 ;
        RECT 0.465000 0.700000 0.535000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.1001 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3471 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.265000 1.040000 0.335000 1.315000 ;
        RECT 0.645000 0.975000 0.715000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.265000 0.085000 0.335000 0.285000 ;
        RECT 0.645000 0.085000 0.715000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085000 0.890000 0.155000 1.250000 ;
      RECT 0.085000 0.820000 0.395000 0.890000 ;
      RECT 0.325000 0.460000 0.395000 0.820000 ;
      RECT 0.085000 0.390000 0.395000 0.460000 ;
      RECT 0.085000 0.150000 0.155000 0.390000 ;
  END
END BUF_X2

MACRO BUF_X32
  CLASS CORE ;
  FOREIGN BUF_X32 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 9.31 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.100000 0.525000 0.170000 0.930000 ;
        RECT 0.100000 0.930000 2.800000 1.000000 ;
        RECT 1.120000 0.560000 1.255000 0.930000 ;
        RECT 1.905000 0.560000 2.040000 0.930000 ;
        RECT 2.665000 0.560000 2.800000 0.930000 ;
    END
    ANTENNAGATEAREA 0.836 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.3672 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1141 LAYER metal1 ;
    ANTENNAGATEAREA 0.836 LAYER metal2 ;
    ANTENNAGATEAREA 0.836 LAYER metal3 ;
    ANTENNAGATEAREA 0.836 LAYER metal4 ;
    ANTENNAGATEAREA 0.836 LAYER metal5 ;
    ANTENNAGATEAREA 0.836 LAYER metal6 ;
    ANTENNAGATEAREA 0.836 LAYER metal7 ;
    ANTENNAGATEAREA 0.836 LAYER metal8 ;
    ANTENNAGATEAREA 0.836 LAYER metal9 ;
    ANTENNAGATEAREA 0.836 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.300000 0.150000 3.370000 0.280000 ;
        RECT 3.300000 0.280000 9.060000 0.420000 ;
        RECT 3.300000 0.420000 3.370000 0.785000 ;
        RECT 3.670000 0.420000 3.740000 0.785000 ;
        RECT 4.050000 0.420000 4.120000 0.785000 ;
        RECT 4.430000 0.420000 4.500000 0.785000 ;
        RECT 4.810000 0.420000 4.880000 0.785000 ;
        RECT 5.190000 0.420000 5.260000 0.785000 ;
        RECT 5.570000 0.420000 5.640000 0.785000 ;
        RECT 5.950000 0.420000 6.020000 0.785000 ;
        RECT 6.330000 0.420000 6.400000 0.785000 ;
        RECT 6.710000 0.420000 6.780000 0.785000 ;
        RECT 7.090000 0.420000 7.160000 0.785000 ;
        RECT 7.470000 0.420000 7.540000 0.785000 ;
        RECT 7.850000 0.420000 7.920000 0.785000 ;
        RECT 8.230000 0.420000 8.300000 0.785000 ;
        RECT 8.610000 0.420000 8.680000 0.785000 ;
        RECT 8.990000 0.420000 9.060000 1.250000 ;
        RECT 3.670000 0.150000 3.740000 0.280000 ;
        RECT 4.050000 0.150000 4.120000 0.280000 ;
        RECT 4.430000 0.150000 4.500000 0.280000 ;
        RECT 4.810000 0.150000 4.880000 0.280000 ;
        RECT 5.190000 0.150000 5.260000 0.280000 ;
        RECT 5.570000 0.150000 5.640000 0.280000 ;
        RECT 5.950000 0.150000 6.020000 0.280000 ;
        RECT 6.330000 0.150000 6.400000 0.280000 ;
        RECT 6.710000 0.150000 6.780000 0.280000 ;
        RECT 7.090000 0.150000 7.160000 0.280000 ;
        RECT 7.470000 0.150000 7.540000 0.280000 ;
        RECT 7.850000 0.150000 7.920000 0.280000 ;
        RECT 8.230000 0.150000 8.300000 0.280000 ;
        RECT 8.610000 0.150000 8.680000 0.280000 ;
        RECT 8.990000 0.150000 9.060000 0.280000 ;
    END
    ANTENNADIFFAREA 2.3617 ;
    ANTENNAPARTIALMETALAREA 1.39335 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 3.7141 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 9.310000 1.485000 ;
        RECT 0.040000 1.065000 0.110000 1.315000 ;
        RECT 0.415000 1.065000 0.485000 1.315000 ;
        RECT 0.795000 1.065000 0.865000 1.315000 ;
        RECT 1.175000 1.065000 1.245000 1.315000 ;
        RECT 1.555000 1.065000 1.625000 1.315000 ;
        RECT 1.935000 1.065000 2.005000 1.315000 ;
        RECT 2.315000 1.065000 2.385000 1.315000 ;
        RECT 2.695000 1.065000 2.765000 1.315000 ;
        RECT 3.080000 1.065000 3.150000 1.315000 ;
        RECT 3.480000 1.065000 3.550000 1.315000 ;
        RECT 3.860000 1.065000 3.930000 1.315000 ;
        RECT 4.240000 1.065000 4.310000 1.315000 ;
        RECT 4.620000 1.065000 4.690000 1.315000 ;
        RECT 5.000000 1.065000 5.070000 1.315000 ;
        RECT 5.380000 1.065000 5.450000 1.315000 ;
        RECT 5.760000 1.065000 5.830000 1.315000 ;
        RECT 6.140000 1.065000 6.210000 1.315000 ;
        RECT 6.520000 1.065000 6.590000 1.315000 ;
        RECT 6.900000 1.065000 6.970000 1.315000 ;
        RECT 7.280000 1.065000 7.350000 1.315000 ;
        RECT 7.660000 1.065000 7.730000 1.315000 ;
        RECT 8.040000 1.065000 8.110000 1.315000 ;
        RECT 8.420000 1.065000 8.490000 1.315000 ;
        RECT 8.800000 1.065000 8.870000 1.315000 ;
        RECT 9.180000 1.065000 9.250000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 9.310000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.360000 ;
        RECT 0.415000 0.085000 0.485000 0.340000 ;
        RECT 0.795000 0.085000 0.865000 0.340000 ;
        RECT 1.175000 0.085000 1.245000 0.340000 ;
        RECT 1.555000 0.085000 1.625000 0.340000 ;
        RECT 1.935000 0.085000 2.005000 0.340000 ;
        RECT 2.315000 0.085000 2.385000 0.340000 ;
        RECT 2.695000 0.085000 2.765000 0.340000 ;
        RECT 3.080000 0.085000 3.150000 0.220000 ;
        RECT 3.480000 0.085000 3.550000 0.200000 ;
        RECT 3.860000 0.085000 3.930000 0.200000 ;
        RECT 4.240000 0.085000 4.310000 0.200000 ;
        RECT 4.620000 0.085000 4.690000 0.200000 ;
        RECT 5.000000 0.085000 5.070000 0.200000 ;
        RECT 5.380000 0.085000 5.450000 0.200000 ;
        RECT 5.760000 0.085000 5.830000 0.200000 ;
        RECT 6.140000 0.085000 6.210000 0.200000 ;
        RECT 6.520000 0.085000 6.590000 0.200000 ;
        RECT 6.900000 0.085000 6.970000 0.200000 ;
        RECT 7.280000 0.085000 7.350000 0.200000 ;
        RECT 7.660000 0.085000 7.730000 0.200000 ;
        RECT 8.040000 0.085000 8.110000 0.200000 ;
        RECT 8.420000 0.085000 8.490000 0.200000 ;
        RECT 8.800000 0.085000 8.870000 0.200000 ;
        RECT 9.180000 0.085000 9.250000 0.200000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 3.165000 0.850000 8.880000 0.920000 ;
      RECT 4.185000 0.560000 4.320000 0.850000 ;
      RECT 5.325000 0.560000 5.460000 0.850000 ;
      RECT 6.465000 0.560000 6.600000 0.850000 ;
      RECT 7.605000 0.560000 7.740000 0.850000 ;
      RECT 8.745000 0.560000 8.880000 0.850000 ;
      RECT 3.165000 0.495000 3.235000 0.850000 ;
      RECT 0.235000 0.405000 3.235000 0.495000 ;
      RECT 0.235000 0.495000 0.305000 0.865000 ;
      RECT 0.615000 0.495000 0.685000 0.865000 ;
      RECT 0.985000 0.495000 1.055000 0.865000 ;
      RECT 1.365000 0.495000 1.435000 0.865000 ;
      RECT 1.745000 0.495000 1.815000 0.865000 ;
      RECT 2.130000 0.495000 2.200000 0.865000 ;
      RECT 2.505000 0.495000 2.575000 0.865000 ;
      RECT 2.885000 0.495000 2.955000 0.865000 ;
      RECT 0.235000 0.150000 0.305000 0.405000 ;
      RECT 0.605000 0.150000 0.675000 0.405000 ;
      RECT 0.985000 0.150000 1.055000 0.405000 ;
      RECT 1.365000 0.150000 1.435000 0.405000 ;
      RECT 1.750000 0.150000 1.820000 0.405000 ;
      RECT 2.130000 0.150000 2.200000 0.405000 ;
      RECT 2.505000 0.150000 2.575000 0.405000 ;
      RECT 2.890000 0.150000 2.960000 0.405000 ;
  END
END BUF_X32

MACRO BUF_X4
  CLASS CORE ;
  FOREIGN BUF_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.170000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615000 0.150000 0.685000 0.560000 ;
        RECT 0.615000 0.560000 1.065000 0.700000 ;
        RECT 0.615000 0.700000 0.685000 1.250000 ;
        RECT 0.995000 0.700000 1.065000 1.250000 ;
        RECT 0.995000 0.150000 1.065000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1974 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6526 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
        RECT 1.175000 0.975000 1.245000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.370000 ;
        RECT 0.415000 0.085000 0.485000 0.370000 ;
        RECT 0.795000 0.085000 0.865000 0.370000 ;
        RECT 1.175000 0.085000 1.245000 0.370000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.660000 0.305000 1.250000 ;
      RECT 0.235000 0.525000 0.550000 0.660000 ;
      RECT 0.235000 0.150000 0.305000 0.525000 ;
  END
END BUF_X4

MACRO BUF_X8
  CLASS CORE ;
  FOREIGN BUF_X8 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.170000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.150000 1.065000 0.560000 ;
        RECT 0.995000 0.560000 2.195000 0.700000 ;
        RECT 0.995000 0.700000 1.065000 1.250000 ;
        RECT 1.365000 0.700000 1.435000 1.250000 ;
        RECT 1.755000 0.700000 1.825000 1.250000 ;
        RECT 2.125000 0.700000 2.195000 1.250000 ;
        RECT 1.365000 0.150000 1.435000 0.560000 ;
        RECT 1.745000 0.150000 1.815000 0.560000 ;
        RECT 2.125000 0.150000 2.195000 0.560000 ;
    END
    ANTENNADIFFAREA 0.5852 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3468 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
        RECT 1.175000 0.975000 1.245000 1.315000 ;
        RECT 1.555000 0.975000 1.625000 1.315000 ;
        RECT 1.935000 0.975000 2.005000 1.315000 ;
        RECT 2.315000 0.975000 2.385000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.415000 0.085000 0.485000 0.425000 ;
        RECT 0.795000 0.085000 0.865000 0.425000 ;
        RECT 1.185000 0.085000 1.255000 0.425000 ;
        RECT 1.555000 0.085000 1.625000 0.425000 ;
        RECT 1.935000 0.085000 2.005000 0.425000 ;
        RECT 2.315000 0.085000 2.385000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.660000 0.305000 1.250000 ;
      RECT 0.235000 0.525000 0.925000 0.660000 ;
      RECT 0.605000 0.660000 0.675000 1.250000 ;
      RECT 0.235000 0.150000 0.305000 0.525000 ;
      RECT 0.605000 0.150000 0.675000 0.525000 ;
  END
END BUF_X8

MACRO CLKBUF_X1
  CLASS CORE ;
  FOREIGN CLKBUF_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.210000 0.700000 ;
    END
    ANTENNAGATEAREA 0.0205 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0845 LAYER metal1 ;
    ANTENNAGATEAREA 0.0205 LAYER metal2 ;
    ANTENNAGATEAREA 0.0205 LAYER metal3 ;
    ANTENNAGATEAREA 0.0205 LAYER metal4 ;
    ANTENNAGATEAREA 0.0205 LAYER metal5 ;
    ANTENNAGATEAREA 0.0205 LAYER metal6 ;
    ANTENNAGATEAREA 0.0205 LAYER metal7 ;
    ANTENNAGATEAREA 0.0205 LAYER metal8 ;
    ANTENNAGATEAREA 0.0205 LAYER metal9 ;
    ANTENNAGATEAREA 0.0205 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.150000 0.510000 1.240000 ;
    END
    ANTENNADIFFAREA 0.086625 ;
    ANTENNAPARTIALMETALAREA 0.0763 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3016 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.570000 1.485000 ;
        RECT 0.245000 0.965000 0.315000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.570000 0.085000 ;
        RECT 0.245000 0.085000 0.315000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.065000 0.900000 0.135000 1.240000 ;
      RECT 0.065000 0.830000 0.370000 0.900000 ;
      RECT 0.300000 0.420000 0.370000 0.830000 ;
      RECT 0.065000 0.350000 0.370000 0.420000 ;
      RECT 0.065000 0.150000 0.135000 0.350000 ;
  END
END CLKBUF_X1

MACRO CLKBUF_X2
  CLASS CORE ;
  FOREIGN CLKBUF_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.190000 0.700000 ;
    END
    ANTENNAGATEAREA 0.04125 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.04125 LAYER metal2 ;
    ANTENNAGATEAREA 0.04125 LAYER metal3 ;
    ANTENNAGATEAREA 0.04125 LAYER metal4 ;
    ANTENNAGATEAREA 0.04125 LAYER metal5 ;
    ANTENNAGATEAREA 0.04125 LAYER metal6 ;
    ANTENNAGATEAREA 0.04125 LAYER metal7 ;
    ANTENNAGATEAREA 0.04125 LAYER metal8 ;
    ANTENNAGATEAREA 0.04125 LAYER metal9 ;
    ANTENNAGATEAREA 0.04125 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.150000 0.510000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1155 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.225000 1.040000 0.295000 1.315000 ;
        RECT 0.605000 0.975000 0.675000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.975000 0.115000 1.250000 ;
      RECT 0.045000 0.905000 0.360000 0.975000 ;
      RECT 0.290000 0.420000 0.360000 0.905000 ;
      RECT 0.045000 0.350000 0.360000 0.420000 ;
      RECT 0.045000 0.150000 0.115000 0.350000 ;
  END
END CLKBUF_X2

MACRO CLKBUF_X3
  CLASS CORE ;
  FOREIGN CLKBUF_X3 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.190000 0.700000 ;
    END
    ANTENNAGATEAREA 0.04125 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.04125 LAYER metal2 ;
    ANTENNAGATEAREA 0.04125 LAYER metal3 ;
    ANTENNAGATEAREA 0.04125 LAYER metal4 ;
    ANTENNAGATEAREA 0.04125 LAYER metal5 ;
    ANTENNAGATEAREA 0.04125 LAYER metal6 ;
    ANTENNAGATEAREA 0.04125 LAYER metal7 ;
    ANTENNAGATEAREA 0.04125 LAYER metal8 ;
    ANTENNAGATEAREA 0.04125 LAYER metal9 ;
    ANTENNAGATEAREA 0.04125 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.180000 0.495000 0.420000 ;
        RECT 0.425000 0.420000 0.865000 0.560000 ;
        RECT 0.425000 0.560000 0.495000 1.175000 ;
        RECT 0.795000 0.560000 0.865000 1.175000 ;
        RECT 0.795000 0.180000 0.865000 0.420000 ;
    END
    ANTENNADIFFAREA 0.202125 ;
    ANTENNAPARTIALMETALAREA 0.1813 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5954 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.225000 0.900000 0.295000 1.315000 ;
        RECT 0.605000 0.900000 0.675000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.235000 ;
        RECT 0.605000 0.085000 0.675000 0.235000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.835000 0.115000 1.175000 ;
      RECT 0.045000 0.765000 0.355000 0.835000 ;
      RECT 0.285000 0.450000 0.355000 0.765000 ;
      RECT 0.045000 0.380000 0.355000 0.450000 ;
      RECT 0.045000 0.180000 0.115000 0.380000 ;
  END
END CLKBUF_X3

MACRO CLKGATETST_X1
  CLASS CORE ;
  FOREIGN CLKGATETST_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.85 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.075000 0.700000 2.220000 0.840000 ;
    END
    ANTENNAGATEAREA 0.0525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.0525 LAYER metal2 ;
    ANTENNAGATEAREA 0.0525 LAYER metal3 ;
    ANTENNAGATEAREA 0.0525 LAYER metal4 ;
    ANTENNAGATEAREA 0.0525 LAYER metal5 ;
    ANTENNAGATEAREA 0.0525 LAYER metal6 ;
    ANTENNAGATEAREA 0.0525 LAYER metal7 ;
    ANTENNAGATEAREA 0.0525 LAYER metal8 ;
    ANTENNAGATEAREA 0.0525 LAYER metal9 ;
    ANTENNAGATEAREA 0.0525 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.700000 0.380000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0182 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.700000 0.185000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SE

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.705000 0.350000 2.790000 1.235000 ;
    END
    ANTENNADIFFAREA 0.086625 ;
    ANTENNAPARTIALMETALAREA 0.075225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2522 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.850000 1.485000 ;
        RECT 2.480000 1.045000 2.615000 1.315000 ;
        RECT 0.385000 1.040000 0.520000 1.315000 ;
        RECT 1.185000 1.010000 1.320000 1.315000 ;
        RECT 1.755000 0.940000 1.825000 1.315000 ;
        RECT 2.135000 0.940000 2.205000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.850000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.420000 ;
        RECT 0.385000 0.085000 0.520000 0.385000 ;
        RECT 1.185000 0.085000 1.320000 0.380000 ;
        RECT 1.750000 0.085000 1.820000 0.420000 ;
        RECT 2.485000 0.085000 2.620000 0.385000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.975000 0.115000 1.235000 ;
      RECT 0.045000 0.905000 0.570000 0.975000 ;
      RECT 0.500000 0.520000 0.570000 0.905000 ;
      RECT 0.235000 0.450000 0.570000 0.520000 ;
      RECT 0.235000 0.285000 0.305000 0.450000 ;
      RECT 0.670000 1.160000 1.120000 1.230000 ;
      RECT 1.050000 0.945000 1.120000 1.160000 ;
      RECT 0.670000 0.220000 0.740000 1.160000 ;
      RECT 1.050000 0.875000 1.475000 0.945000 ;
      RECT 0.670000 0.150000 1.015000 0.220000 ;
      RECT 1.405000 0.945000 1.475000 1.235000 ;
      RECT 0.945000 0.220000 1.015000 0.445000 ;
      RECT 0.945000 0.445000 1.475000 0.515000 ;
      RECT 1.405000 0.285000 1.475000 0.445000 ;
      RECT 0.805000 0.805000 0.875000 1.095000 ;
      RECT 0.805000 0.735000 1.555000 0.805000 ;
      RECT 0.805000 0.285000 0.875000 0.735000 ;
      RECT 1.565000 0.930000 1.690000 1.205000 ;
      RECT 1.620000 0.655000 1.690000 0.930000 ;
      RECT 1.105000 0.585000 1.690000 0.655000 ;
      RECT 1.565000 0.285000 1.635000 0.585000 ;
      RECT 1.935000 0.220000 2.005000 1.210000 ;
      RECT 1.935000 0.150000 2.070000 0.220000 ;
      RECT 2.330000 0.660000 2.400000 1.005000 ;
      RECT 2.330000 0.595000 2.640000 0.660000 ;
      RECT 2.140000 0.525000 2.640000 0.595000 ;
      RECT 2.140000 0.285000 2.210000 0.525000 ;
  END
END CLKGATETST_X1

MACRO CLKGATETST_X2
  CLASS CORE ;
  FOREIGN CLKGATETST_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.04 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.180000 0.525000 2.250000 0.850000 ;
        RECT 2.180000 0.850000 2.825000 0.920000 ;
        RECT 2.720000 0.525000 2.825000 0.850000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.102025 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3549 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.560000 0.375000 0.725000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.020625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0754 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.560000 0.545000 0.725000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.017325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0702 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SE

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.520000 0.150000 2.600000 0.785000 ;
    END
    ANTENNADIFFAREA 0.1155 ;
    ANTENNAPARTIALMETALAREA 0.0508 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1859 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.040000 1.485000 ;
        RECT 1.830000 1.240000 1.965000 1.315000 ;
        RECT 2.275000 1.240000 2.410000 1.315000 ;
        RECT 2.675000 1.240000 2.810000 1.315000 ;
        RECT 0.730000 1.115000 0.865000 1.315000 ;
        RECT 0.225000 0.940000 0.295000 1.315000 ;
        RECT 1.515000 0.910000 1.585000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.040000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.285000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
        RECT 1.450000 0.085000 1.520000 0.405000 ;
        RECT 1.765000 0.085000 1.900000 0.185000 ;
        RECT 2.325000 0.085000 2.395000 0.195000 ;
        RECT 2.700000 0.085000 2.770000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.610000 0.545000 0.680000 0.885000 ;
      RECT 0.610000 0.480000 0.870000 0.545000 ;
      RECT 0.425000 0.410000 0.870000 0.480000 ;
      RECT 0.425000 0.150000 0.495000 0.410000 ;
      RECT 0.045000 0.875000 0.115000 1.125000 ;
      RECT 0.045000 0.805000 0.480000 0.875000 ;
      RECT 0.410000 0.875000 0.480000 0.950000 ;
      RECT 0.045000 0.150000 0.115000 0.805000 ;
      RECT 0.410000 0.950000 1.015000 1.020000 ;
      RECT 0.945000 0.745000 1.015000 0.950000 ;
      RECT 0.945000 0.610000 1.080000 0.745000 ;
      RECT 0.945000 0.220000 1.015000 0.610000 ;
      RECT 0.945000 0.150000 1.285000 0.220000 ;
      RECT 1.145000 0.660000 1.215000 1.030000 ;
      RECT 1.145000 0.525000 1.630000 0.660000 ;
      RECT 1.145000 0.420000 1.215000 0.525000 ;
      RECT 1.080000 0.285000 1.215000 0.420000 ;
      RECT 1.380000 0.760000 1.775000 0.830000 ;
      RECT 1.705000 0.350000 1.775000 0.760000 ;
      RECT 1.610000 0.280000 1.775000 0.350000 ;
      RECT 2.045000 0.460000 2.115000 0.925000 ;
      RECT 2.045000 0.390000 2.450000 0.460000 ;
      RECT 2.170000 0.325000 2.450000 0.390000 ;
      RECT 2.170000 0.150000 2.240000 0.325000 ;
      RECT 1.680000 1.150000 1.750000 1.245000 ;
      RECT 1.680000 1.080000 2.965000 1.150000 ;
      RECT 2.895000 1.150000 2.965000 1.240000 ;
      RECT 2.895000 0.150000 2.965000 1.080000 ;
  END
END CLKGATETST_X2

MACRO CLKGATETST_X4
  CLASS CORE ;
  FOREIGN CLKGATETST_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.210000 0.525000 2.280000 0.770000 ;
        RECT 2.210000 0.770000 2.850000 0.850000 ;
        RECT 2.720000 0.525000 2.850000 0.770000 ;
    END
    ANTENNAGATEAREA 0.13075 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1002 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3146 LAYER metal1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal2 ;
    ANTENNAGATEAREA 0.13075 LAYER metal3 ;
    ANTENNAGATEAREA 0.13075 LAYER metal4 ;
    ANTENNAGATEAREA 0.13075 LAYER metal5 ;
    ANTENNAGATEAREA 0.13075 LAYER metal6 ;
    ANTENNAGATEAREA 0.13075 LAYER metal7 ;
    ANTENNAGATEAREA 0.13075 LAYER metal8 ;
    ANTENNAGATEAREA 0.13075 LAYER metal9 ;
    ANTENNAGATEAREA 0.13075 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.560000 0.380000 0.775000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02795 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0897 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.560000 0.185000 0.775000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.026875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0884 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SE

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.085000 0.180000 3.155000 0.420000 ;
        RECT 3.085000 0.420000 3.525000 0.560000 ;
        RECT 3.085000 0.560000 3.155000 0.925000 ;
        RECT 3.455000 0.560000 3.525000 0.925000 ;
        RECT 3.455000 0.180000 3.525000 0.420000 ;
    END
    ANTENNADIFFAREA 0.231 ;
    ANTENNAPARTIALMETALAREA 0.1463 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4654 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.800000 1.485000 ;
        RECT 2.130000 1.205000 2.200000 1.315000 ;
        RECT 2.505000 1.200000 2.575000 1.315000 ;
        RECT 2.885000 1.200000 2.955000 1.315000 ;
        RECT 1.490000 1.165000 1.625000 1.315000 ;
        RECT 0.755000 1.130000 0.825000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 3.265000 0.975000 3.335000 1.315000 ;
        RECT 3.645000 0.975000 3.715000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.800000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.285000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.755000 0.085000 0.825000 0.195000 ;
        RECT 1.530000 0.085000 1.600000 0.285000 ;
        RECT 2.125000 0.085000 2.195000 0.285000 ;
        RECT 2.885000 0.085000 2.955000 0.200000 ;
        RECT 3.265000 0.085000 3.335000 0.200000 ;
        RECT 3.645000 0.085000 3.715000 0.200000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.910000 0.115000 1.250000 ;
      RECT 0.045000 0.840000 0.910000 0.910000 ;
      RECT 0.840000 0.485000 0.910000 0.840000 ;
      RECT 0.235000 0.415000 0.910000 0.485000 ;
      RECT 0.235000 0.150000 0.335000 0.415000 ;
      RECT 0.575000 1.045000 0.645000 1.250000 ;
      RECT 0.575000 0.975000 1.065000 1.045000 ;
      RECT 0.975000 0.460000 1.065000 0.975000 ;
      RECT 0.975000 0.390000 1.325000 0.460000 ;
      RECT 0.975000 0.330000 1.045000 0.390000 ;
      RECT 0.575000 0.260000 1.045000 0.330000 ;
      RECT 0.575000 0.150000 0.645000 0.260000 ;
      RECT 1.405000 0.725000 1.780000 0.795000 ;
      RECT 1.710000 0.150000 1.780000 0.725000 ;
      RECT 1.265000 0.865000 1.990000 0.935000 ;
      RECT 1.265000 0.795000 1.335000 0.865000 ;
      RECT 1.920000 0.150000 1.990000 0.865000 ;
      RECT 1.130000 1.100000 1.205000 1.250000 ;
      RECT 1.130000 1.030000 2.125000 1.100000 ;
      RECT 1.130000 0.660000 1.200000 1.030000 ;
      RECT 2.055000 0.460000 2.125000 1.030000 ;
      RECT 1.130000 0.525000 1.645000 0.660000 ;
      RECT 2.055000 0.390000 2.495000 0.460000 ;
      RECT 1.390000 0.255000 1.460000 0.525000 ;
      RECT 2.425000 0.460000 2.495000 0.660000 ;
      RECT 1.110000 0.185000 1.460000 0.255000 ;
      RECT 2.290000 0.930000 3.015000 1.000000 ;
      RECT 2.945000 0.420000 3.015000 0.930000 ;
      RECT 2.655000 0.350000 3.015000 0.420000 ;
      RECT 2.655000 0.255000 2.725000 0.350000 ;
      RECT 2.480000 0.185000 2.725000 0.255000 ;
  END
END CLKGATETST_X4

MACRO CLKGATETST_X8
  CLASS CORE ;
  FOREIGN CLKGATETST_X8 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 5.51 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.385000 0.525000 2.455000 0.845000 ;
        RECT 2.385000 0.845000 3.925000 0.915000 ;
        RECT 3.100000 0.630000 3.170000 0.845000 ;
        RECT 3.855000 0.630000 3.925000 0.845000 ;
        RECT 3.035000 0.560000 3.170000 0.630000 ;
        RECT 3.765000 0.560000 3.925000 0.630000 ;
    END
    ANTENNAGATEAREA 0.23525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.18095 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6903 LAYER metal1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal2 ;
    ANTENNAGATEAREA 0.23525 LAYER metal3 ;
    ANTENNAGATEAREA 0.23525 LAYER metal4 ;
    ANTENNAGATEAREA 0.23525 LAYER metal5 ;
    ANTENNAGATEAREA 0.23525 LAYER metal6 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ;
    ANTENNAGATEAREA 0.23525 LAYER metal8 ;
    ANTENNAGATEAREA 0.23525 LAYER metal9 ;
    ANTENNAGATEAREA 0.23525 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.330000 0.700000 0.510000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0252 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.700000 0.250000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0266 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END SE

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.075000 0.975000 4.190000 1.250000 ;
        RECT 4.120000 0.700000 4.190000 0.975000 ;
        RECT 4.120000 0.560000 5.275000 0.700000 ;
        RECT 4.445000 0.700000 4.515000 1.250000 ;
        RECT 4.825000 0.700000 4.895000 1.250000 ;
        RECT 5.205000 0.700000 5.275000 1.250000 ;
        RECT 4.120000 0.285000 4.190000 0.560000 ;
        RECT 4.445000 0.150000 4.515000 0.560000 ;
        RECT 4.825000 0.150000 4.895000 0.560000 ;
        RECT 5.205000 0.150000 5.275000 0.560000 ;
        RECT 4.075000 0.150000 4.190000 0.285000 ;
    END
    ANTENNADIFFAREA 0.462 ;
    ANTENNAPARTIALMETALAREA 0.44895 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3585 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 5.510000 1.485000 ;
        RECT 0.750000 1.240000 0.885000 1.315000 ;
        RECT 0.410000 1.215000 0.545000 1.315000 ;
        RECT 1.535000 1.100000 1.670000 1.315000 ;
        RECT 1.915000 1.100000 2.050000 1.315000 ;
        RECT 2.365000 1.060000 2.435000 1.315000 ;
        RECT 2.705000 1.010000 2.840000 1.315000 ;
        RECT 3.085000 1.010000 3.220000 1.315000 ;
        RECT 3.465000 1.010000 3.600000 1.315000 ;
        RECT 3.845000 1.010000 3.980000 1.315000 ;
        RECT 4.260000 0.975000 4.330000 1.315000 ;
        RECT 4.635000 0.975000 4.705000 1.315000 ;
        RECT 5.015000 0.975000 5.085000 1.315000 ;
        RECT 5.395000 0.975000 5.465000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 5.510000 0.085000 ;
        RECT 0.065000 0.085000 0.135000 0.285000 ;
        RECT 0.440000 0.085000 0.510000 0.285000 ;
        RECT 0.750000 0.085000 0.885000 0.175000 ;
        RECT 1.575000 0.085000 1.645000 0.265000 ;
        RECT 1.950000 0.085000 2.020000 0.425000 ;
        RECT 2.330000 0.085000 2.465000 0.160000 ;
        RECT 3.085000 0.085000 3.220000 0.160000 ;
        RECT 3.845000 0.085000 3.980000 0.250000 ;
        RECT 4.255000 0.085000 4.325000 0.285000 ;
        RECT 4.635000 0.085000 4.705000 0.285000 ;
        RECT 5.015000 0.085000 5.085000 0.285000 ;
        RECT 5.395000 0.085000 5.465000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.070000 0.975000 0.140000 1.250000 ;
      RECT 0.070000 0.905000 0.950000 0.975000 ;
      RECT 0.870000 0.490000 0.950000 0.905000 ;
      RECT 0.260000 0.420000 0.950000 0.490000 ;
      RECT 0.260000 0.150000 0.330000 0.420000 ;
      RECT 0.565000 1.065000 1.085000 1.135000 ;
      RECT 1.015000 0.495000 1.085000 1.065000 ;
      RECT 1.015000 0.425000 1.370000 0.495000 ;
      RECT 1.015000 0.320000 1.085000 0.425000 ;
      RECT 0.600000 0.250000 1.085000 0.320000 ;
      RECT 0.600000 0.150000 0.670000 0.250000 ;
      RECT 1.450000 0.695000 1.885000 0.765000 ;
      RECT 1.815000 0.390000 1.885000 0.695000 ;
      RECT 1.730000 0.185000 1.885000 0.390000 ;
      RECT 1.315000 0.830000 2.170000 0.900000 ;
      RECT 1.315000 0.715000 1.385000 0.830000 ;
      RECT 2.100000 0.195000 2.170000 0.830000 ;
      RECT 1.160000 1.035000 1.230000 1.185000 ;
      RECT 1.160000 0.965000 2.305000 1.035000 ;
      RECT 1.160000 0.630000 1.230000 0.965000 ;
      RECT 2.235000 0.360000 2.305000 0.965000 ;
      RECT 1.160000 0.560000 1.750000 0.630000 ;
      RECT 2.235000 0.290000 3.440000 0.360000 ;
      RECT 1.435000 0.250000 1.505000 0.560000 ;
      RECT 2.575000 0.360000 2.645000 0.560000 ;
      RECT 3.370000 0.360000 3.440000 0.555000 ;
      RECT 1.155000 0.180000 1.505000 0.250000 ;
      RECT 2.575000 0.560000 2.735000 0.630000 ;
      RECT 3.370000 0.555000 3.520000 0.625000 ;
      RECT 2.520000 0.710000 3.030000 0.780000 ;
      RECT 2.900000 0.495000 2.970000 0.710000 ;
      RECT 2.710000 0.425000 3.305000 0.495000 ;
      RECT 3.235000 0.495000 3.305000 0.705000 ;
      RECT 3.235000 0.705000 3.700000 0.710000 ;
      RECT 3.235000 0.710000 3.790000 0.780000 ;
      RECT 3.630000 0.485000 3.700000 0.705000 ;
      RECT 3.630000 0.350000 4.055000 0.485000 ;
      RECT 3.630000 0.230000 3.700000 0.350000 ;
      RECT 3.470000 0.160000 3.700000 0.230000 ;
  END
END CLKGATETST_X8

MACRO CLKGATE_X1
  CLASS CORE ;
  FOREIGN CLKGATE_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.540000 0.420000 1.895000 0.560000 ;
    END
    ANTENNAGATEAREA 0.0525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0497 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1287 LAYER metal1 ;
    ANTENNAGATEAREA 0.0525 LAYER metal2 ;
    ANTENNAGATEAREA 0.0525 LAYER metal3 ;
    ANTENNAGATEAREA 0.0525 LAYER metal4 ;
    ANTENNAGATEAREA 0.0525 LAYER metal5 ;
    ANTENNAGATEAREA 0.0525 LAYER metal6 ;
    ANTENNAGATEAREA 0.0525 LAYER metal7 ;
    ANTENNAGATEAREA 0.0525 LAYER metal8 ;
    ANTENNAGATEAREA 0.0525 LAYER metal9 ;
    ANTENNAGATEAREA 0.0525 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.910000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0897 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.310000 0.175000 2.410000 1.090000 ;
    END
    ANTENNADIFFAREA 0.086625 ;
    ANTENNAPARTIALMETALAREA 0.0915 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2639 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.225000 0.955000 0.295000 1.315000 ;
        RECT 2.030000 0.915000 2.100000 1.315000 ;
        RECT 0.955000 0.900000 1.090000 1.315000 ;
        RECT 1.585000 0.890000 1.655000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.320000 ;
        RECT 0.985000 0.085000 1.055000 0.320000 ;
        RECT 1.585000 0.085000 1.655000 0.195000 ;
        RECT 2.120000 0.085000 2.190000 0.225000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.040000 0.520000 0.110000 1.040000 ;
      RECT 0.040000 0.450000 0.440000 0.520000 ;
      RECT 0.040000 0.265000 0.110000 0.450000 ;
      RECT 0.510000 0.980000 0.715000 1.050000 ;
      RECT 0.510000 0.725000 0.580000 0.980000 ;
      RECT 0.175000 0.590000 0.580000 0.725000 ;
      RECT 0.510000 0.290000 0.580000 0.590000 ;
      RECT 0.510000 0.220000 0.710000 0.290000 ;
      RECT 1.175000 0.835000 1.245000 1.050000 ;
      RECT 0.695000 0.765000 1.245000 0.835000 ;
      RECT 0.695000 0.460000 0.765000 0.765000 ;
      RECT 0.695000 0.390000 1.245000 0.460000 ;
      RECT 1.175000 0.270000 1.245000 0.390000 ;
      RECT 1.405000 0.660000 1.475000 1.090000 ;
      RECT 1.145000 0.525000 1.475000 0.660000 ;
      RECT 1.405000 0.195000 1.475000 0.525000 ;
      RECT 1.785000 0.835000 1.855000 1.090000 ;
      RECT 1.785000 0.765000 2.245000 0.835000 ;
      RECT 2.175000 0.420000 2.245000 0.765000 ;
      RECT 1.970000 0.350000 2.245000 0.420000 ;
      RECT 1.970000 0.185000 2.040000 0.350000 ;
  END
END CLKGATE_X1

MACRO CLKGATE_X2
  CLASS CORE ;
  FOREIGN CLKGATE_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.580000 0.420000 1.650000 0.660000 ;
    END
    ANTENNAGATEAREA 0.0785 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0168 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.0785 LAYER metal2 ;
    ANTENNAGATEAREA 0.0785 LAYER metal3 ;
    ANTENNAGATEAREA 0.0785 LAYER metal4 ;
    ANTENNAGATEAREA 0.0785 LAYER metal5 ;
    ANTENNAGATEAREA 0.0785 LAYER metal6 ;
    ANTENNAGATEAREA 0.0785 LAYER metal7 ;
    ANTENNAGATEAREA 0.0785 LAYER metal8 ;
    ANTENNAGATEAREA 0.0785 LAYER metal9 ;
    ANTENNAGATEAREA 0.0785 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.340000 0.420000 0.510000 0.590000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0289 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0884 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.320000 0.185000 2.410000 1.215000 ;
    END
    ANTENNADIFFAREA 0.1155 ;
    ANTENNAPARTIALMETALAREA 0.0927 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2912 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.660000 1.485000 ;
        RECT 0.985000 0.980000 1.055000 1.315000 ;
        RECT 0.225000 0.940000 0.295000 1.315000 ;
        RECT 2.095000 0.940000 2.165000 1.315000 ;
        RECT 2.505000 0.940000 2.575000 1.315000 ;
        RECT 1.725000 0.890000 1.795000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.660000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.320000 ;
        RECT 0.955000 0.085000 1.090000 0.285000 ;
        RECT 1.565000 0.085000 1.635000 0.235000 ;
        RECT 2.095000 0.085000 2.165000 0.220000 ;
        RECT 2.505000 0.085000 2.575000 0.220000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.605000 0.725000 0.675000 1.115000 ;
      RECT 0.175000 0.655000 0.675000 0.725000 ;
      RECT 0.175000 0.525000 0.245000 0.655000 ;
      RECT 0.605000 0.200000 0.675000 0.655000 ;
      RECT 1.255000 0.720000 1.325000 1.115000 ;
      RECT 0.740000 0.650000 1.325000 0.720000 ;
      RECT 0.740000 0.585000 0.990000 0.650000 ;
      RECT 0.920000 0.420000 0.990000 0.585000 ;
      RECT 0.920000 0.350000 1.280000 0.420000 ;
      RECT 1.420000 0.560000 1.490000 0.975000 ;
      RECT 1.065000 0.490000 1.490000 0.560000 ;
      RECT 1.385000 0.185000 1.455000 0.490000 ;
      RECT 0.360000 1.180000 0.920000 1.250000 ;
      RECT 0.360000 0.875000 0.430000 1.180000 ;
      RECT 0.850000 0.860000 0.920000 1.180000 ;
      RECT 0.040000 0.805000 0.430000 0.875000 ;
      RECT 0.850000 0.790000 1.190000 0.860000 ;
      RECT 0.040000 0.875000 0.110000 1.170000 ;
      RECT 0.040000 0.295000 0.110000 0.805000 ;
      RECT 1.120000 0.860000 1.190000 1.180000 ;
      RECT 1.120000 1.180000 1.640000 1.250000 ;
      RECT 1.570000 0.825000 1.640000 1.180000 ;
      RECT 1.570000 0.755000 1.785000 0.825000 ;
      RECT 1.715000 0.630000 1.785000 0.755000 ;
      RECT 1.715000 0.560000 2.095000 0.630000 ;
      RECT 1.915000 0.875000 1.985000 1.215000 ;
      RECT 1.915000 0.805000 2.255000 0.875000 ;
      RECT 2.185000 0.460000 2.255000 0.805000 ;
      RECT 1.725000 0.390000 2.255000 0.460000 ;
      RECT 1.725000 0.185000 1.795000 0.390000 ;
  END
END CLKGATE_X2

MACRO CLKGATE_X4
  CLASS CORE ;
  FOREIGN CLKGATE_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.535000 0.390000 1.965000 0.460000 ;
        RECT 1.535000 0.460000 1.650000 0.700000 ;
        RECT 1.895000 0.460000 1.965000 0.660000 ;
    END
    ANTENNAGATEAREA 0.13075 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0717 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2444 LAYER metal1 ;
    ANTENNAGATEAREA 0.13075 LAYER metal2 ;
    ANTENNAGATEAREA 0.13075 LAYER metal3 ;
    ANTENNAGATEAREA 0.13075 LAYER metal4 ;
    ANTENNAGATEAREA 0.13075 LAYER metal5 ;
    ANTENNAGATEAREA 0.13075 LAYER metal6 ;
    ANTENNAGATEAREA 0.13075 LAYER metal7 ;
    ANTENNAGATEAREA 0.13075 LAYER metal8 ;
    ANTENNAGATEAREA 0.13075 LAYER metal9 ;
    ANTENNAGATEAREA 0.13075 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.350000 0.420000 0.510000 0.630000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0336 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0962 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END E

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.555000 0.150000 2.625000 0.420000 ;
        RECT 2.555000 0.420000 2.995000 0.560000 ;
        RECT 2.555000 0.560000 2.625000 1.240000 ;
        RECT 2.925000 0.560000 2.995000 1.240000 ;
        RECT 2.925000 0.150000 2.995000 0.420000 ;
    END
    ANTENNADIFFAREA 0.231 ;
    ANTENNAPARTIALMETALAREA 0.1946 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6448 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.230000 1.485000 ;
        RECT 1.570000 1.240000 1.705000 1.315000 ;
        RECT 1.975000 1.065000 2.045000 1.315000 ;
        RECT 2.355000 1.065000 2.425000 1.315000 ;
        RECT 0.235000 0.965000 0.305000 1.315000 ;
        RECT 0.995000 0.965000 1.065000 1.315000 ;
        RECT 2.735000 0.965000 2.805000 1.315000 ;
        RECT 3.115000 0.965000 3.185000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.230000 0.085000 ;
        RECT 0.235000 0.085000 0.305000 0.320000 ;
        RECT 0.995000 0.085000 1.065000 0.320000 ;
        RECT 1.580000 0.085000 1.650000 0.285000 ;
        RECT 2.325000 0.085000 2.460000 0.185000 ;
        RECT 2.735000 0.085000 2.805000 0.215000 ;
        RECT 3.115000 0.085000 3.185000 0.215000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.615000 0.765000 0.685000 1.095000 ;
      RECT 0.185000 0.695000 0.685000 0.765000 ;
      RECT 0.185000 0.525000 0.255000 0.695000 ;
      RECT 0.615000 0.200000 0.685000 0.695000 ;
      RECT 1.265000 0.765000 1.335000 0.870000 ;
      RECT 1.055000 0.695000 1.335000 0.765000 ;
      RECT 1.055000 0.460000 1.125000 0.695000 ;
      RECT 0.750000 0.390000 1.255000 0.460000 ;
      RECT 0.750000 0.460000 0.820000 0.660000 ;
      RECT 1.185000 0.300000 1.255000 0.390000 ;
      RECT 1.400000 0.630000 1.470000 1.040000 ;
      RECT 1.190000 0.560000 1.470000 0.630000 ;
      RECT 1.400000 0.150000 1.470000 0.560000 ;
      RECT 0.370000 1.165000 0.885000 1.235000 ;
      RECT 0.370000 0.900000 0.440000 1.165000 ;
      RECT 0.815000 0.900000 0.885000 1.165000 ;
      RECT 0.050000 0.830000 0.440000 0.900000 ;
      RECT 0.815000 0.830000 1.200000 0.900000 ;
      RECT 0.050000 0.900000 0.120000 1.240000 ;
      RECT 0.050000 0.150000 0.120000 0.830000 ;
      RECT 1.130000 0.900000 1.200000 1.105000 ;
      RECT 0.920000 0.560000 0.990000 0.830000 ;
      RECT 1.130000 1.105000 1.640000 1.175000 ;
      RECT 1.570000 0.835000 1.640000 1.105000 ;
      RECT 1.570000 0.765000 2.320000 0.835000 ;
      RECT 1.715000 0.525000 1.785000 0.765000 ;
      RECT 2.250000 0.525000 2.320000 0.765000 ;
      RECT 1.790000 0.975000 1.860000 1.240000 ;
      RECT 1.790000 0.905000 2.490000 0.975000 ;
      RECT 2.165000 0.975000 2.235000 1.240000 ;
      RECT 2.420000 0.325000 2.490000 0.905000 ;
      RECT 1.950000 0.255000 2.490000 0.325000 ;
  END
END CLKGATE_X4

MACRO CLKGATE_X8
  CLASS CORE ;
  FOREIGN CLKGATE_X8 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.625000 0.860000 2.935000 0.930000 ;
        RECT 2.130000 0.525000 2.220000 0.860000 ;
        RECT 2.865000 0.525000 2.935000 0.860000 ;
    END
    ANTENNAGATEAREA 0.23525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1453 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.533 LAYER metal1 ;
    ANTENNAGATEAREA 0.23525 LAYER metal2 ;
    ANTENNAGATEAREA 0.23525 LAYER metal3 ;
    ANTENNAGATEAREA 0.23525 LAYER metal4 ;
    ANTENNAGATEAREA 0.23525 LAYER metal5 ;
    ANTENNAGATEAREA 0.23525 LAYER metal6 ;
    ANTENNAGATEAREA 0.23525 LAYER metal7 ;
    ANTENNAGATEAREA 0.23525 LAYER metal8 ;
    ANTENNAGATEAREA 0.23525 LAYER metal9 ;
    ANTENNAGATEAREA 0.23525 LAYER metal10 ;
  END CK

  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.345000 0.560000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END E

  PIN GCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.485000 0.150000 3.555000 0.420000 ;
        RECT 3.485000 0.420000 4.685000 0.560000 ;
        RECT 3.485000 0.560000 3.555000 1.235000 ;
        RECT 3.855000 0.560000 3.925000 1.235000 ;
        RECT 4.235000 0.560000 4.305000 1.235000 ;
        RECT 4.615000 0.560000 4.685000 1.235000 ;
        RECT 3.855000 0.150000 3.925000 0.420000 ;
        RECT 4.235000 0.150000 4.305000 0.420000 ;
        RECT 4.615000 0.150000 4.685000 0.420000 ;
    END
    ANTENNADIFFAREA 0.462 ;
    ANTENNAPARTIALMETALAREA 0.4326 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3312 LAYER metal1 ;
  END GCK

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.940000 1.485000 ;
        RECT 2.120000 1.205000 2.190000 1.315000 ;
        RECT 2.500000 1.205000 2.570000 1.315000 ;
        RECT 2.880000 1.205000 2.950000 1.315000 ;
        RECT 1.355000 1.175000 1.490000 1.315000 ;
        RECT 1.725000 1.065000 1.795000 1.315000 ;
        RECT 1.005000 0.995000 1.075000 1.315000 ;
        RECT 0.230000 0.960000 0.300000 1.315000 ;
        RECT 3.275000 0.960000 3.345000 1.315000 ;
        RECT 3.665000 0.960000 3.735000 1.315000 ;
        RECT 4.045000 0.960000 4.115000 1.315000 ;
        RECT 4.425000 0.960000 4.495000 1.315000 ;
        RECT 4.805000 0.960000 4.875000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.940000 0.085000 ;
        RECT 0.200000 0.085000 0.335000 0.250000 ;
        RECT 1.005000 0.085000 1.075000 0.285000 ;
        RECT 1.355000 0.085000 1.490000 0.160000 ;
        RECT 1.715000 0.085000 1.850000 0.160000 ;
        RECT 2.470000 0.085000 2.605000 0.160000 ;
        RECT 3.245000 0.085000 3.380000 0.160000 ;
        RECT 3.670000 0.085000 3.740000 0.285000 ;
        RECT 4.045000 0.085000 4.115000 0.285000 ;
        RECT 4.425000 0.085000 4.495000 0.285000 ;
        RECT 4.805000 0.085000 4.875000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.460000 0.115000 1.235000 ;
      RECT 0.045000 0.390000 0.800000 0.460000 ;
      RECT 0.575000 0.460000 0.645000 0.870000 ;
      RECT 0.045000 0.150000 0.115000 0.390000 ;
      RECT 0.585000 1.010000 0.805000 1.080000 ;
      RECT 0.735000 0.660000 0.805000 1.010000 ;
      RECT 0.735000 0.525000 1.140000 0.660000 ;
      RECT 0.865000 0.250000 0.935000 0.525000 ;
      RECT 0.585000 0.180000 0.935000 0.250000 ;
      RECT 0.440000 1.150000 0.940000 1.220000 ;
      RECT 0.870000 0.930000 0.940000 1.150000 ;
      RECT 0.440000 0.835000 0.510000 1.150000 ;
      RECT 0.870000 0.860000 1.560000 0.930000 ;
      RECT 0.180000 0.765000 0.510000 0.835000 ;
      RECT 1.490000 0.930000 1.560000 1.005000 ;
      RECT 1.490000 0.500000 1.560000 0.860000 ;
      RECT 0.180000 0.605000 0.250000 0.765000 ;
      RECT 1.490000 1.005000 1.645000 1.075000 ;
      RECT 1.490000 0.430000 1.645000 0.500000 ;
      RECT 0.870000 0.725000 1.275000 0.795000 ;
      RECT 1.205000 0.325000 1.275000 0.725000 ;
      RECT 1.205000 0.255000 3.225000 0.325000 ;
      RECT 1.825000 0.325000 1.895000 0.660000 ;
      RECT 2.500000 0.325000 2.570000 0.660000 ;
      RECT 3.155000 0.325000 3.225000 0.660000 ;
      RECT 1.205000 0.150000 1.275000 0.255000 ;
      RECT 1.905000 1.065000 2.040000 1.200000 ;
      RECT 1.905000 0.995000 3.140000 1.065000 ;
      RECT 2.280000 1.065000 2.415000 1.200000 ;
      RECT 2.660000 1.065000 2.795000 1.200000 ;
      RECT 3.070000 1.065000 3.140000 1.235000 ;
      RECT 3.070000 0.795000 3.140000 0.995000 ;
      RECT 3.005000 0.725000 3.420000 0.795000 ;
      RECT 3.350000 0.525000 3.420000 0.725000 ;
      RECT 3.005000 0.460000 3.075000 0.725000 ;
      RECT 2.670000 0.390000 3.075000 0.460000 ;
      RECT 2.670000 0.460000 2.740000 0.725000 ;
      RECT 2.310000 0.725000 2.740000 0.795000 ;
      RECT 2.310000 0.460000 2.380000 0.725000 ;
      RECT 2.095000 0.390000 2.380000 0.460000 ;
  END
END CLKGATE_X8

MACRO DFFRS_X1
  CLASS CORE ;
  FOREIGN DFFRS_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.56 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.120000 0.585000 4.310000 0.840000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.04845 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1157 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.200000 0.700000 1.345000 0.840000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END RN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.800000 0.700000 0.890000 0.840000 ;
    END
    ANTENNAGATEAREA 0.0615 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0126 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0598 LAYER metal1 ;
    ANTENNAGATEAREA 0.0615 LAYER metal2 ;
    ANTENNAGATEAREA 0.0615 LAYER metal3 ;
    ANTENNAGATEAREA 0.0615 LAYER metal4 ;
    ANTENNAGATEAREA 0.0615 LAYER metal5 ;
    ANTENNAGATEAREA 0.0615 LAYER metal6 ;
    ANTENNAGATEAREA 0.0615 LAYER metal7 ;
    ANTENNAGATEAREA 0.0615 LAYER metal8 ;
    ANTENNAGATEAREA 0.0615 LAYER metal9 ;
    ANTENNAGATEAREA 0.0615 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.240000 0.280000 4.385000 0.495000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.031175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0936 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.400000 0.510000 0.875000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.03325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1417 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.185000 0.130000 1.075000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0623 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2496 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.560000 1.485000 ;
        RECT 0.215000 1.100000 0.350000 1.315000 ;
        RECT 0.560000 1.095000 0.695000 1.315000 ;
        RECT 0.965000 1.065000 1.035000 1.315000 ;
        RECT 3.325000 1.030000 3.460000 1.315000 ;
        RECT 1.655000 0.990000 1.790000 1.315000 ;
        RECT 1.345000 0.925000 1.415000 1.315000 ;
        RECT 4.255000 0.915000 4.325000 1.315000 ;
        RECT 2.415000 0.890000 2.550000 1.315000 ;
        RECT 2.795000 0.835000 2.930000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.560000 0.085000 ;
        RECT 0.215000 0.085000 0.350000 0.200000 ;
        RECT 0.935000 0.085000 1.070000 0.285000 ;
        RECT 1.470000 0.085000 1.605000 0.285000 ;
        RECT 2.415000 0.085000 2.550000 0.285000 ;
        RECT 3.135000 0.085000 3.270000 0.285000 ;
        RECT 4.225000 0.085000 4.360000 0.160000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200000 0.960000 0.880000 1.030000 ;
      RECT 0.200000 0.335000 0.270000 0.960000 ;
      RECT 0.200000 0.265000 0.695000 0.335000 ;
      RECT 0.955000 0.925000 1.260000 0.995000 ;
      RECT 0.955000 0.625000 1.025000 0.925000 ;
      RECT 0.595000 0.555000 1.025000 0.625000 ;
      RECT 0.950000 0.425000 1.025000 0.555000 ;
      RECT 0.950000 0.350000 1.900000 0.425000 ;
      RECT 1.505000 0.925000 1.575000 1.075000 ;
      RECT 1.505000 0.855000 1.945000 0.925000 ;
      RECT 1.875000 0.925000 1.945000 1.075000 ;
      RECT 2.065000 0.630000 2.135000 1.085000 ;
      RECT 1.090000 0.495000 2.135000 0.630000 ;
      RECT 2.065000 0.185000 2.135000 0.495000 ;
      RECT 2.635000 0.825000 2.705000 1.070000 ;
      RECT 2.345000 0.755000 2.705000 0.825000 ;
      RECT 2.345000 0.555000 2.415000 0.755000 ;
      RECT 2.345000 0.485000 3.545000 0.555000 ;
      RECT 2.825000 0.300000 2.895000 0.485000 ;
      RECT 3.175000 0.965000 3.245000 1.115000 ;
      RECT 3.175000 0.895000 3.615000 0.965000 ;
      RECT 3.545000 0.965000 3.615000 1.115000 ;
      RECT 3.850000 0.690000 3.920000 1.115000 ;
      RECT 2.500000 0.620000 3.920000 0.690000 ;
      RECT 3.760000 0.285000 3.830000 0.620000 ;
      RECT 1.955000 1.165000 2.275000 1.235000 ;
      RECT 2.205000 0.420000 2.275000 1.165000 ;
      RECT 2.205000 0.350000 2.760000 0.420000 ;
      RECT 2.690000 0.235000 2.760000 0.350000 ;
      RECT 2.690000 0.165000 3.050000 0.235000 ;
      RECT 2.980000 0.235000 3.050000 0.350000 ;
      RECT 2.980000 0.350000 3.690000 0.420000 ;
      RECT 3.620000 0.420000 3.690000 0.460000 ;
      RECT 3.620000 0.220000 3.690000 0.350000 ;
      RECT 3.620000 0.150000 4.055000 0.220000 ;
      RECT 3.985000 0.220000 4.055000 1.180000 ;
      RECT 3.680000 1.180000 4.055000 1.250000 ;
      RECT 3.680000 0.830000 3.750000 1.180000 ;
      RECT 3.020000 0.760000 3.750000 0.830000 ;
      RECT 3.020000 0.830000 3.090000 1.070000 ;
      RECT 4.450000 0.185000 4.520000 1.250000 ;
  END
END DFFRS_X1

MACRO DFFRS_X2
  CLASS CORE ;
  FOREIGN DFFRS_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.94 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.485000 0.280000 4.690000 0.460000 ;
        RECT 4.485000 0.460000 4.555000 0.575000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.04495 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.390000 0.545000 1.460000 0.700000 ;
    END
    ANTENNAGATEAREA 0.04875 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01085 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAGATEAREA 0.04875 LAYER metal2 ;
    ANTENNAGATEAREA 0.04875 LAYER metal3 ;
    ANTENNAGATEAREA 0.04875 LAYER metal4 ;
    ANTENNAGATEAREA 0.04875 LAYER metal5 ;
    ANTENNAGATEAREA 0.04875 LAYER metal6 ;
    ANTENNAGATEAREA 0.04875 LAYER metal7 ;
    ANTENNAGATEAREA 0.04875 LAYER metal8 ;
    ANTENNAGATEAREA 0.04875 LAYER metal9 ;
    ANTENNAGATEAREA 0.04875 LAYER metal10 ;
  END RN

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.200000 0.545000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.075 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01085 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0585 LAYER metal1 ;
    ANTENNAGATEAREA 0.075 LAYER metal2 ;
    ANTENNAGATEAREA 0.075 LAYER metal3 ;
    ANTENNAGATEAREA 0.075 LAYER metal4 ;
    ANTENNAGATEAREA 0.075 LAYER metal5 ;
    ANTENNAGATEAREA 0.075 LAYER metal6 ;
    ANTENNAGATEAREA 0.075 LAYER metal7 ;
    ANTENNAGATEAREA 0.075 LAYER metal8 ;
    ANTENNAGATEAREA 0.075 LAYER metal9 ;
    ANTENNAGATEAREA 0.075 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 4.620000 0.540000 4.720000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.016 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.625000 0.400000 0.700000 0.965000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.042375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1664 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.240000 0.200000 0.320000 0.965000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0612 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2197 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.940000 1.485000 ;
        RECT 0.425000 1.205000 0.495000 1.315000 ;
        RECT 0.875000 1.205000 0.945000 1.315000 ;
        RECT 1.335000 1.080000 1.405000 1.315000 ;
        RECT 3.695000 1.030000 3.830000 1.315000 ;
        RECT 2.055000 0.955000 2.125000 1.315000 ;
        RECT 2.815000 0.955000 2.885000 1.315000 ;
        RECT 0.050000 0.925000 0.120000 1.315000 ;
        RECT 1.715000 0.895000 1.785000 1.315000 ;
        RECT 3.195000 0.765000 3.265000 1.315000 ;
        RECT 4.590000 0.765000 4.660000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.940000 0.085000 ;
        RECT 0.050000 0.085000 0.120000 0.415000 ;
        RECT 0.425000 0.085000 0.495000 0.200000 ;
        RECT 0.805000 0.085000 0.875000 0.200000 ;
        RECT 1.335000 0.085000 1.405000 0.320000 ;
        RECT 1.870000 0.085000 1.940000 0.320000 ;
        RECT 2.785000 0.085000 2.920000 0.285000 ;
        RECT 3.505000 0.085000 3.640000 0.285000 ;
        RECT 4.560000 0.085000 4.695000 0.215000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.490000 1.035000 1.225000 1.105000 ;
      RECT 0.490000 0.660000 0.560000 1.035000 ;
      RECT 0.385000 0.525000 0.560000 0.660000 ;
      RECT 0.490000 0.335000 0.560000 0.525000 ;
      RECT 0.490000 0.265000 1.065000 0.335000 ;
      RECT 1.065000 0.845000 1.630000 0.915000 ;
      RECT 1.065000 0.660000 1.135000 0.845000 ;
      RECT 0.840000 0.525000 1.135000 0.660000 ;
      RECT 1.065000 0.480000 1.135000 0.525000 ;
      RECT 1.065000 0.410000 2.270000 0.480000 ;
      RECT 1.715000 0.205000 1.785000 0.410000 ;
      RECT 1.875000 0.890000 1.945000 1.075000 ;
      RECT 1.875000 0.820000 2.315000 0.890000 ;
      RECT 2.245000 0.890000 2.315000 1.075000 ;
      RECT 2.425000 0.650000 2.505000 1.075000 ;
      RECT 1.580000 0.580000 2.505000 0.650000 ;
      RECT 2.425000 0.200000 2.505000 0.580000 ;
      RECT 3.005000 0.825000 3.075000 1.040000 ;
      RECT 2.760000 0.755000 3.075000 0.825000 ;
      RECT 2.760000 0.555000 2.830000 0.755000 ;
      RECT 2.760000 0.485000 3.915000 0.555000 ;
      RECT 3.195000 0.320000 3.265000 0.485000 ;
      RECT 3.545000 0.965000 3.615000 1.115000 ;
      RECT 3.545000 0.895000 3.985000 0.965000 ;
      RECT 3.915000 0.965000 3.985000 1.115000 ;
      RECT 4.185000 0.690000 4.255000 1.115000 ;
      RECT 2.895000 0.620000 4.255000 0.690000 ;
      RECT 4.130000 0.285000 4.200000 0.620000 ;
      RECT 2.325000 1.140000 2.640000 1.210000 ;
      RECT 2.570000 0.420000 2.640000 1.140000 ;
      RECT 2.570000 0.350000 3.130000 0.420000 ;
      RECT 3.060000 0.255000 3.130000 0.350000 ;
      RECT 3.060000 0.185000 3.420000 0.255000 ;
      RECT 3.350000 0.255000 3.420000 0.350000 ;
      RECT 3.350000 0.350000 4.055000 0.420000 ;
      RECT 3.985000 0.420000 4.055000 0.460000 ;
      RECT 3.985000 0.220000 4.055000 0.350000 ;
      RECT 3.985000 0.150000 4.390000 0.220000 ;
      RECT 4.320000 0.220000 4.390000 1.180000 ;
      RECT 4.050000 1.180000 4.390000 1.250000 ;
      RECT 4.050000 0.830000 4.120000 1.180000 ;
      RECT 3.390000 0.760000 4.120000 0.830000 ;
      RECT 3.390000 0.830000 3.460000 1.040000 ;
      RECT 4.785000 0.250000 4.855000 1.240000 ;
  END
END DFFRS_X2

MACRO DFFR_X1
  CLASS CORE ;
  FOREIGN DFFR_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.600000 0.560000 0.720000 0.745000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0222 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.495000 1.165000 1.885000 1.235000 ;
        RECT 1.815000 1.000000 1.885000 1.165000 ;
        RECT 1.815000 0.930000 2.175000 1.000000 ;
        RECT 2.105000 1.000000 2.175000 1.180000 ;
        RECT 2.105000 1.180000 2.525000 1.250000 ;
        RECT 2.455000 0.710000 2.525000 1.180000 ;
        RECT 2.455000 0.640000 2.890000 0.710000 ;
        RECT 2.455000 0.560000 2.600000 0.640000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.181 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6682 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END RN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.175000 0.420000 0.320000 0.560000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0203 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.660000 0.185000 3.740000 1.250000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0852 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2977 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.285000 0.400000 3.360000 1.250000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.06375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2405 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.800000 1.485000 ;
        RECT 0.230000 1.065000 0.300000 1.315000 ;
        RECT 1.950000 1.065000 2.020000 1.315000 ;
        RECT 3.080000 1.065000 3.150000 1.315000 ;
        RECT 1.295000 1.030000 1.430000 1.315000 ;
        RECT 0.575000 1.015000 0.645000 1.315000 ;
        RECT 2.700000 0.980000 2.770000 1.315000 ;
        RECT 3.465000 0.975000 3.535000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.800000 0.085000 ;
        RECT 0.230000 0.085000 0.300000 0.320000 ;
        RECT 0.575000 0.085000 0.645000 0.320000 ;
        RECT 1.515000 0.085000 1.585000 0.410000 ;
        RECT 1.895000 0.085000 2.030000 0.285000 ;
        RECT 2.700000 0.085000 2.770000 0.320000 ;
        RECT 3.465000 0.085000 3.535000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.040000 0.835000 0.110000 1.250000 ;
      RECT 0.040000 0.700000 0.355000 0.835000 ;
      RECT 0.040000 0.185000 0.110000 0.700000 ;
      RECT 1.495000 1.025000 1.630000 1.095000 ;
      RECT 1.495000 0.965000 1.565000 1.025000 ;
      RECT 1.135000 0.895000 1.565000 0.965000 ;
      RECT 1.135000 0.965000 1.205000 1.125000 ;
      RECT 0.955000 0.695000 1.025000 1.125000 ;
      RECT 0.955000 0.625000 1.895000 0.695000 ;
      RECT 0.955000 0.290000 1.025000 0.625000 ;
      RECT 1.985000 0.555000 2.120000 0.670000 ;
      RECT 1.090000 0.485000 2.120000 0.555000 ;
      RECT 1.090000 0.220000 1.160000 0.485000 ;
      RECT 0.820000 0.150000 1.160000 0.220000 ;
      RECT 0.820000 0.220000 0.890000 0.425000 ;
      RECT 0.420000 0.425000 0.890000 0.495000 ;
      RECT 0.420000 0.495000 0.490000 1.250000 ;
      RECT 0.820000 0.495000 0.890000 0.785000 ;
      RECT 0.420000 0.185000 0.490000 0.425000 ;
      RECT 1.680000 0.830000 1.750000 0.960000 ;
      RECT 1.190000 0.760000 2.255000 0.830000 ;
      RECT 2.185000 0.420000 2.255000 0.760000 ;
      RECT 1.690000 0.350000 2.255000 0.420000 ;
      RECT 1.690000 0.185000 1.760000 0.350000 ;
      RECT 2.320000 0.495000 2.390000 1.115000 ;
      RECT 2.320000 0.425000 3.050000 0.495000 ;
      RECT 2.980000 0.495000 3.050000 0.660000 ;
      RECT 2.320000 0.185000 2.390000 0.425000 ;
      RECT 2.890000 0.880000 2.960000 1.250000 ;
      RECT 2.590000 0.810000 3.185000 0.880000 ;
      RECT 3.115000 0.335000 3.185000 0.810000 ;
      RECT 3.050000 0.265000 3.595000 0.335000 ;
      RECT 3.525000 0.335000 3.595000 0.660000 ;
  END
END DFFR_X1

MACRO DFFR_X2
  CLASS CORE ;
  FOREIGN DFFR_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 4.18 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.520000 0.740000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0198 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0754 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.515000 1.165000 1.905000 1.235000 ;
        RECT 1.835000 1.035000 1.905000 1.165000 ;
        RECT 1.835000 0.965000 2.240000 1.035000 ;
        RECT 2.170000 1.035000 2.240000 1.150000 ;
        RECT 2.170000 1.150000 2.590000 1.220000 ;
        RECT 2.520000 0.700000 2.590000 1.150000 ;
        RECT 2.520000 0.560000 2.905000 0.700000 ;
    END
    ANTENNAGATEAREA 0.06125 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1876 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6331 LAYER metal1 ;
    ANTENNAGATEAREA 0.06125 LAYER metal2 ;
    ANTENNAGATEAREA 0.06125 LAYER metal3 ;
    ANTENNAGATEAREA 0.06125 LAYER metal4 ;
    ANTENNAGATEAREA 0.06125 LAYER metal5 ;
    ANTENNAGATEAREA 0.06125 LAYER metal6 ;
    ANTENNAGATEAREA 0.06125 LAYER metal7 ;
    ANTENNAGATEAREA 0.06125 LAYER metal8 ;
    ANTENNAGATEAREA 0.06125 LAYER metal9 ;
    ANTENNAGATEAREA 0.06125 LAYER metal10 ;
  END RN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.195000 0.420000 0.320000 0.560000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.860000 0.185000 3.935000 1.080000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.067125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2522 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.410000 0.645000 3.550000 0.785000 ;
        RECT 3.480000 0.185000 3.550000 0.645000 ;
    END
    ANTENNADIFFAREA 0.1904 ;
    ANTENNAPARTIALMETALAREA 0.0518 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1924 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 4.180000 1.485000 ;
        RECT 1.970000 1.100000 2.105000 1.315000 ;
        RECT 3.190000 1.065000 3.260000 1.315000 ;
        RECT 3.670000 1.065000 3.740000 1.315000 ;
        RECT 4.050000 1.065000 4.120000 1.315000 ;
        RECT 1.315000 1.030000 1.450000 1.315000 ;
        RECT 0.590000 1.015000 0.660000 1.315000 ;
        RECT 2.725000 1.000000 2.860000 1.315000 ;
        RECT 0.245000 0.945000 0.315000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 4.180000 0.085000 ;
        RECT 0.245000 0.085000 0.315000 0.320000 ;
        RECT 0.590000 0.085000 0.660000 0.320000 ;
        RECT 1.535000 0.085000 1.605000 0.410000 ;
        RECT 1.900000 0.085000 2.035000 0.285000 ;
        RECT 2.690000 0.085000 2.760000 0.320000 ;
        RECT 3.295000 0.085000 3.365000 0.195000 ;
        RECT 3.670000 0.085000 3.740000 0.335000 ;
        RECT 4.050000 0.085000 4.120000 0.335000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 0.790000 0.130000 1.220000 ;
      RECT 0.060000 0.655000 0.375000 0.790000 ;
      RECT 0.060000 0.185000 0.130000 0.655000 ;
      RECT 1.515000 1.025000 1.650000 1.095000 ;
      RECT 1.515000 0.965000 1.585000 1.025000 ;
      RECT 1.155000 0.895000 1.585000 0.965000 ;
      RECT 1.155000 0.965000 1.225000 1.125000 ;
      RECT 0.970000 0.695000 1.040000 1.125000 ;
      RECT 0.970000 0.625000 1.925000 0.695000 ;
      RECT 1.850000 0.695000 1.925000 0.765000 ;
      RECT 0.970000 0.290000 1.040000 0.625000 ;
      RECT 2.055000 0.555000 2.125000 0.705000 ;
      RECT 1.105000 0.485000 2.125000 0.555000 ;
      RECT 1.105000 0.220000 1.175000 0.485000 ;
      RECT 0.830000 0.150000 1.175000 0.220000 ;
      RECT 0.830000 0.220000 0.900000 0.385000 ;
      RECT 0.440000 0.385000 0.900000 0.455000 ;
      RECT 0.440000 0.455000 0.510000 0.980000 ;
      RECT 0.830000 0.455000 0.900000 0.820000 ;
      RECT 0.440000 0.185000 0.510000 0.385000 ;
      RECT 1.700000 0.900000 1.770000 0.960000 ;
      RECT 1.700000 0.830000 2.260000 0.900000 ;
      RECT 1.235000 0.760000 1.770000 0.830000 ;
      RECT 2.190000 0.420000 2.260000 0.830000 ;
      RECT 1.750000 0.350000 2.260000 0.420000 ;
      RECT 1.750000 0.185000 1.820000 0.350000 ;
      RECT 2.375000 0.455000 2.445000 1.085000 ;
      RECT 2.375000 0.385000 2.950000 0.455000 ;
      RECT 2.880000 0.335000 2.950000 0.385000 ;
      RECT 2.375000 0.285000 2.445000 0.385000 ;
      RECT 2.880000 0.265000 3.310000 0.335000 ;
      RECT 2.285000 0.215000 2.445000 0.285000 ;
      RECT 3.240000 0.335000 3.310000 0.660000 ;
      RECT 2.970000 0.920000 3.040000 1.220000 ;
      RECT 2.655000 0.850000 3.790000 0.920000 ;
      RECT 2.655000 0.765000 2.725000 0.850000 ;
      RECT 3.720000 0.525000 3.790000 0.850000 ;
      RECT 3.070000 0.400000 3.140000 0.850000 ;
  END
END DFFR_X2

MACRO DFFS_X1
  CLASS CORE ;
  FOREIGN DFFS_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.340000 0.560000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0238 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.625000 0.700000 2.790000 0.840000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.705000 0.590000 1.840000 0.725000 ;
        RECT 1.770000 0.725000 1.840000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.026275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1001 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.575000 0.185000 3.645000 0.560000 ;
        RECT 3.575000 0.560000 3.740000 0.700000 ;
        RECT 3.575000 0.700000 3.645000 1.160000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.08155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2964 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.195000 0.185000 3.265000 0.560000 ;
        RECT 3.195000 0.560000 3.360000 0.700000 ;
        RECT 3.195000 0.700000 3.265000 0.925000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0651 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2353 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.800000 1.485000 ;
        RECT 3.380000 1.205000 3.450000 1.315000 ;
        RECT 2.480000 1.065000 2.615000 1.315000 ;
        RECT 2.855000 1.005000 2.925000 1.315000 ;
        RECT 1.015000 0.940000 1.085000 1.315000 ;
        RECT 1.755000 0.905000 1.825000 1.315000 ;
        RECT 0.225000 0.900000 0.295000 1.315000 ;
        RECT 1.410000 0.885000 1.480000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.800000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.320000 ;
        RECT 1.040000 0.085000 1.110000 0.320000 ;
        RECT 1.750000 0.085000 1.820000 0.375000 ;
        RECT 2.670000 0.085000 2.805000 0.340000 ;
        RECT 3.385000 0.085000 3.455000 0.460000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.040000 0.835000 0.110000 1.160000 ;
      RECT 0.040000 0.765000 0.570000 0.835000 ;
      RECT 0.040000 0.185000 0.110000 0.765000 ;
      RECT 0.590000 0.975000 0.865000 1.045000 ;
      RECT 0.795000 0.615000 0.865000 0.975000 ;
      RECT 0.770000 0.545000 1.350000 0.615000 ;
      RECT 1.280000 0.615000 1.350000 0.685000 ;
      RECT 0.770000 0.355000 0.840000 0.545000 ;
      RECT 0.590000 0.285000 0.840000 0.355000 ;
      RECT 1.220000 0.820000 1.290000 1.090000 ;
      RECT 0.940000 0.750000 1.485000 0.820000 ;
      RECT 0.940000 0.685000 1.010000 0.750000 ;
      RECT 1.415000 0.285000 1.485000 0.750000 ;
      RECT 1.570000 0.815000 1.670000 1.090000 ;
      RECT 1.570000 0.510000 1.640000 0.815000 ;
      RECT 1.570000 0.440000 2.040000 0.510000 ;
      RECT 1.970000 0.510000 2.040000 0.665000 ;
      RECT 1.570000 0.220000 1.640000 0.440000 ;
      RECT 1.970000 0.220000 2.040000 0.440000 ;
      RECT 1.970000 0.665000 2.095000 0.800000 ;
      RECT 1.280000 0.150000 1.640000 0.220000 ;
      RECT 1.970000 0.150000 2.320000 0.220000 ;
      RECT 1.280000 0.220000 1.350000 0.385000 ;
      RECT 0.905000 0.385000 1.350000 0.455000 ;
      RECT 0.905000 0.220000 0.975000 0.385000 ;
      RECT 0.445000 0.150000 0.975000 0.220000 ;
      RECT 0.445000 0.220000 0.515000 0.420000 ;
      RECT 0.175000 0.420000 0.705000 0.490000 ;
      RECT 0.175000 0.490000 0.245000 0.685000 ;
      RECT 0.635000 0.490000 0.705000 0.720000 ;
      RECT 0.635000 0.720000 0.730000 0.855000 ;
      RECT 2.330000 1.000000 2.400000 1.150000 ;
      RECT 2.330000 0.930000 2.770000 1.000000 ;
      RECT 2.700000 1.000000 2.770000 1.150000 ;
      RECT 2.105000 1.045000 2.240000 1.115000 ;
      RECT 2.170000 0.630000 2.240000 1.045000 ;
      RECT 2.170000 0.560000 2.925000 0.630000 ;
      RECT 2.170000 0.360000 2.240000 0.560000 ;
      RECT 2.105000 0.290000 2.240000 0.360000 ;
      RECT 3.010000 0.995000 3.505000 1.065000 ;
      RECT 3.435000 0.525000 3.505000 0.995000 ;
      RECT 3.010000 0.490000 3.080000 0.995000 ;
      RECT 2.375000 0.420000 3.080000 0.490000 ;
      RECT 2.905000 0.185000 2.975000 0.420000 ;
  END
END DFFS_X1

MACRO DFFS_X2
  CLASS CORE ;
  FOREIGN DFFS_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.99 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.350000 0.560000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0224 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.675000 0.560000 2.790000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03525 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0161 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0663 LAYER metal1 ;
    ANTENNAGATEAREA 0.03525 LAYER metal2 ;
    ANTENNAGATEAREA 0.03525 LAYER metal3 ;
    ANTENNAGATEAREA 0.03525 LAYER metal4 ;
    ANTENNAGATEAREA 0.03525 LAYER metal5 ;
    ANTENNAGATEAREA 0.03525 LAYER metal6 ;
    ANTENNAGATEAREA 0.03525 LAYER metal7 ;
    ANTENNAGATEAREA 0.03525 LAYER metal8 ;
    ANTENNAGATEAREA 0.03525 LAYER metal9 ;
    ANTENNAGATEAREA 0.03525 LAYER metal10 ;
  END SN

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.750000 0.590000 1.840000 0.840000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0225 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0884 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.100000 0.400000 3.170000 0.925000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.03675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1547 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.480000 0.400000 3.550000 0.925000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.03675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1547 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.990000 1.485000 ;
        RECT 2.910000 1.205000 2.980000 1.315000 ;
        RECT 3.285000 1.205000 3.355000 1.315000 ;
        RECT 3.660000 1.205000 3.730000 1.315000 ;
        RECT 2.530000 1.065000 2.665000 1.315000 ;
        RECT 0.235000 0.940000 0.305000 1.315000 ;
        RECT 1.080000 0.940000 1.150000 1.315000 ;
        RECT 1.460000 0.940000 1.530000 1.315000 ;
        RECT 1.805000 0.940000 1.875000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.990000 0.085000 ;
        RECT 0.235000 0.085000 0.305000 0.320000 ;
        RECT 1.090000 0.085000 1.160000 0.370000 ;
        RECT 1.800000 0.085000 1.870000 0.320000 ;
        RECT 2.720000 0.085000 2.855000 0.340000 ;
        RECT 3.280000 0.085000 3.350000 0.195000 ;
        RECT 3.660000 0.085000 3.730000 0.195000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.050000 0.835000 0.120000 1.215000 ;
      RECT 0.050000 0.765000 0.585000 0.835000 ;
      RECT 0.050000 0.185000 0.120000 0.765000 ;
      RECT 0.585000 0.975000 0.890000 1.045000 ;
      RECT 0.820000 0.705000 0.890000 0.975000 ;
      RECT 0.820000 0.570000 1.400000 0.705000 ;
      RECT 0.820000 0.355000 0.890000 0.570000 ;
      RECT 0.590000 0.285000 0.890000 0.355000 ;
      RECT 0.965000 0.770000 1.535000 0.840000 ;
      RECT 1.465000 0.285000 1.535000 0.770000 ;
      RECT 1.615000 0.940000 1.720000 1.075000 ;
      RECT 1.615000 0.525000 1.685000 0.940000 ;
      RECT 1.615000 0.455000 2.090000 0.525000 ;
      RECT 2.020000 0.525000 2.090000 0.665000 ;
      RECT 1.615000 0.220000 1.685000 0.455000 ;
      RECT 2.020000 0.220000 2.090000 0.455000 ;
      RECT 2.020000 0.665000 2.145000 0.800000 ;
      RECT 1.225000 0.150000 1.685000 0.220000 ;
      RECT 2.020000 0.150000 2.395000 0.220000 ;
      RECT 1.225000 0.220000 1.295000 0.435000 ;
      RECT 0.955000 0.435000 1.295000 0.505000 ;
      RECT 0.955000 0.220000 1.025000 0.435000 ;
      RECT 0.455000 0.150000 1.025000 0.220000 ;
      RECT 0.455000 0.220000 0.525000 0.425000 ;
      RECT 0.190000 0.425000 0.720000 0.495000 ;
      RECT 0.190000 0.495000 0.260000 0.695000 ;
      RECT 0.650000 0.495000 0.720000 0.735000 ;
      RECT 0.650000 0.735000 0.755000 0.870000 ;
      RECT 2.380000 1.000000 2.450000 1.150000 ;
      RECT 2.380000 0.930000 2.820000 1.000000 ;
      RECT 2.750000 1.000000 2.820000 1.150000 ;
      RECT 2.155000 1.045000 2.290000 1.115000 ;
      RECT 2.220000 0.475000 2.290000 1.045000 ;
      RECT 2.220000 0.405000 3.035000 0.475000 ;
      RECT 2.220000 0.360000 2.290000 0.405000 ;
      RECT 2.965000 0.335000 3.035000 0.405000 ;
      RECT 2.155000 0.290000 2.290000 0.360000 ;
      RECT 2.965000 0.265000 3.685000 0.335000 ;
      RECT 3.615000 0.335000 3.685000 0.660000 ;
      RECT 3.850000 1.060000 3.920000 1.215000 ;
      RECT 2.920000 0.990000 3.920000 1.060000 ;
      RECT 2.920000 0.865000 2.990000 0.990000 ;
      RECT 3.235000 0.525000 3.305000 0.990000 ;
      RECT 3.850000 0.260000 3.920000 0.990000 ;
      RECT 2.450000 0.795000 2.990000 0.865000 ;
  END
END DFFS_X2

MACRO DFF_X1
  CLASS CORE ;
  FOREIGN DFF_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.810000 0.530000 0.970000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0272 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.560000 0.530000 1.670000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0187 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.100000 0.260000 3.170000 1.130000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0609 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2444 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.720000 0.260000 2.790000 0.785000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.03675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1547 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.230000 1.485000 ;
        RECT 2.345000 1.100000 2.480000 1.315000 ;
        RECT 1.005000 1.080000 1.075000 1.315000 ;
        RECT 2.905000 0.985000 2.975000 1.315000 ;
        RECT 0.240000 0.980000 0.310000 1.315000 ;
        RECT 1.610000 0.900000 1.680000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.230000 0.085000 ;
        RECT 0.240000 0.085000 0.310000 0.405000 ;
        RECT 0.975000 0.085000 1.110000 0.300000 ;
        RECT 1.610000 0.085000 1.680000 0.360000 ;
        RECT 2.345000 0.085000 2.480000 0.370000 ;
        RECT 2.905000 0.085000 2.975000 0.460000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 0.745000 0.130000 1.130000 ;
      RECT 0.060000 0.610000 0.570000 0.745000 ;
      RECT 0.060000 0.270000 0.130000 0.610000 ;
      RECT 0.635000 0.835000 0.705000 1.115000 ;
      RECT 0.635000 0.765000 1.190000 0.835000 ;
      RECT 1.120000 0.530000 1.190000 0.765000 ;
      RECT 0.635000 0.285000 0.705000 0.765000 ;
      RECT 1.275000 0.440000 1.345000 0.995000 ;
      RECT 0.785000 0.370000 1.345000 0.440000 ;
      RECT 1.200000 0.270000 1.270000 0.370000 ;
      RECT 0.785000 0.220000 0.855000 0.370000 ;
      RECT 0.380000 0.150000 0.855000 0.220000 ;
      RECT 0.380000 0.220000 0.450000 0.545000 ;
      RECT 0.485000 1.180000 0.940000 1.250000 ;
      RECT 0.870000 1.015000 0.940000 1.180000 ;
      RECT 0.870000 0.945000 1.210000 1.015000 ;
      RECT 1.140000 1.015000 1.210000 1.180000 ;
      RECT 1.140000 1.180000 1.495000 1.250000 ;
      RECT 1.425000 0.835000 1.495000 1.180000 ;
      RECT 1.425000 0.765000 1.925000 0.835000 ;
      RECT 1.425000 0.225000 1.495000 0.765000 ;
      RECT 1.855000 0.220000 1.925000 0.765000 ;
      RECT 1.855000 0.150000 2.205000 0.220000 ;
      RECT 2.000000 0.660000 2.070000 1.200000 ;
      RECT 2.000000 0.525000 2.505000 0.660000 ;
      RECT 2.000000 0.285000 2.070000 0.525000 ;
      RECT 2.570000 0.920000 2.640000 1.115000 ;
      RECT 2.570000 0.850000 3.035000 0.920000 ;
      RECT 2.570000 0.800000 2.640000 0.850000 ;
      RECT 2.965000 0.525000 3.035000 0.850000 ;
      RECT 2.265000 0.730000 2.640000 0.800000 ;
      RECT 2.570000 0.225000 2.640000 0.730000 ;
  END
END DFF_X1

MACRO DFF_X2
  CLASS CORE ;
  FOREIGN DFF_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.61 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.940000 0.560000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.570000 0.560000 1.650000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0112 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0572 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END CK

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.290000 0.250000 3.360000 1.115000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.06055 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2431 LAYER metal1 ;
  END Q

  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.910000 0.250000 2.980000 0.925000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.04725 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1937 LAYER metal1 ;
  END QN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.610000 1.485000 ;
        RECT 2.730000 1.205000 2.800000 1.315000 ;
        RECT 3.105000 1.205000 3.175000 1.315000 ;
        RECT 1.015000 1.080000 1.085000 1.315000 ;
        RECT 0.255000 0.965000 0.325000 1.315000 ;
        RECT 1.620000 0.900000 1.690000 1.315000 ;
        RECT 2.350000 0.875000 2.485000 1.315000 ;
        RECT 3.485000 0.840000 3.555000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.610000 0.085000 ;
        RECT 0.255000 0.085000 0.325000 0.385000 ;
        RECT 0.985000 0.085000 1.120000 0.215000 ;
        RECT 1.620000 0.085000 1.690000 0.385000 ;
        RECT 2.350000 0.085000 2.485000 0.450000 ;
        RECT 2.730000 0.085000 2.800000 0.460000 ;
        RECT 3.105000 0.085000 3.175000 0.460000 ;
        RECT 3.485000 0.085000 3.555000 0.460000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.075000 0.835000 0.145000 1.055000 ;
      RECT 0.075000 0.765000 0.625000 0.835000 ;
      RECT 0.555000 0.565000 0.625000 0.765000 ;
      RECT 0.075000 0.325000 0.145000 0.765000 ;
      RECT 0.610000 1.000000 0.760000 1.070000 ;
      RECT 0.690000 0.835000 0.760000 1.000000 ;
      RECT 0.690000 0.765000 1.215000 0.835000 ;
      RECT 1.145000 0.565000 1.215000 0.765000 ;
      RECT 0.690000 0.355000 0.760000 0.765000 ;
      RECT 0.610000 0.285000 0.760000 0.355000 ;
      RECT 1.285000 0.355000 1.355000 1.115000 ;
      RECT 0.825000 0.285000 1.355000 0.355000 ;
      RECT 0.825000 0.220000 0.895000 0.285000 ;
      RECT 0.390000 0.150000 0.895000 0.220000 ;
      RECT 0.390000 0.220000 0.460000 0.700000 ;
      RECT 0.500000 1.180000 0.935000 1.250000 ;
      RECT 0.865000 1.015000 0.935000 1.180000 ;
      RECT 0.865000 0.945000 1.220000 1.015000 ;
      RECT 1.150000 1.015000 1.220000 1.180000 ;
      RECT 1.150000 1.180000 1.505000 1.250000 ;
      RECT 1.435000 0.835000 1.505000 1.180000 ;
      RECT 1.435000 0.765000 1.945000 0.835000 ;
      RECT 1.875000 0.285000 1.945000 0.765000 ;
      RECT 1.435000 0.250000 1.505000 0.765000 ;
      RECT 1.875000 0.215000 2.215000 0.285000 ;
      RECT 2.010000 0.660000 2.080000 0.975000 ;
      RECT 2.010000 0.525000 2.510000 0.660000 ;
      RECT 2.010000 0.350000 2.080000 0.525000 ;
      RECT 2.575000 1.045000 3.215000 1.115000 ;
      RECT 2.575000 0.805000 2.645000 1.045000 ;
      RECT 3.145000 0.525000 3.215000 1.045000 ;
      RECT 2.245000 0.735000 2.645000 0.805000 ;
      RECT 2.575000 0.200000 2.645000 0.735000 ;
  END
END DFF_X2

MACRO DLH_X1
  CLASS CORE ;
  FOREIGN DLH_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.9 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.950000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.200000 0.525000 0.320000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0767 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END G

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.185000 0.510000 0.785000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.042 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1742 LAYER metal1 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.900000 1.485000 ;
        RECT 1.595000 1.025000 1.665000 1.315000 ;
        RECT 0.250000 0.985000 0.320000 1.315000 ;
        RECT 0.845000 0.965000 0.915000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.900000 0.085000 ;
        RECT 0.250000 0.085000 0.320000 0.320000 ;
        RECT 0.805000 0.085000 0.940000 0.285000 ;
        RECT 1.595000 0.085000 1.665000 0.445000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.505000 1.180000 0.780000 1.250000 ;
      RECT 0.505000 0.920000 0.575000 1.180000 ;
      RECT 0.065000 0.850000 0.575000 0.920000 ;
      RECT 0.065000 0.920000 0.135000 1.240000 ;
      RECT 0.065000 0.185000 0.135000 0.850000 ;
      RECT 1.025000 1.180000 1.430000 1.250000 ;
      RECT 1.025000 0.835000 1.095000 1.180000 ;
      RECT 0.650000 0.765000 1.215000 0.835000 ;
      RECT 0.650000 0.835000 0.720000 1.115000 ;
      RECT 1.145000 0.560000 1.215000 0.765000 ;
      RECT 0.650000 0.185000 0.720000 0.765000 ;
      RECT 1.145000 0.490000 1.280000 0.560000 ;
      RECT 1.190000 1.045000 1.415000 1.115000 ;
      RECT 1.345000 0.795000 1.415000 1.045000 ;
      RECT 1.345000 0.660000 1.725000 0.795000 ;
      RECT 1.345000 0.420000 1.415000 0.660000 ;
      RECT 0.785000 0.350000 1.415000 0.420000 ;
      RECT 0.785000 0.420000 0.855000 0.660000 ;
      RECT 1.790000 0.595000 1.860000 1.160000 ;
      RECT 1.485000 0.525000 1.860000 0.595000 ;
      RECT 1.790000 0.320000 1.860000 0.525000 ;
  END
END DLH_X1

MACRO DLH_X2
  CLASS CORE ;
  FOREIGN DLH_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.135000 0.525000 1.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.03475 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.023625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.03475 LAYER metal2 ;
    ANTENNAGATEAREA 0.03475 LAYER metal3 ;
    ANTENNAGATEAREA 0.03475 LAYER metal4 ;
    ANTENNAGATEAREA 0.03475 LAYER metal5 ;
    ANTENNAGATEAREA 0.03475 LAYER metal6 ;
    ANTENNAGATEAREA 0.03475 LAYER metal7 ;
    ANTENNAGATEAREA 0.03475 LAYER metal8 ;
    ANTENNAGATEAREA 0.03475 LAYER metal9 ;
    ANTENNAGATEAREA 0.03475 LAYER metal10 ;
  END D

  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.180000 0.525000 0.320000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0819 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END G

  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.185000 0.510000 0.785000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.042 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1742 LAYER metal1 ;
  END Q

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 1.780000 1.080000 1.850000 1.315000 ;
        RECT 0.240000 1.055000 0.310000 1.315000 ;
        RECT 1.030000 1.040000 1.100000 1.315000 ;
        RECT 0.620000 1.000000 0.690000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.240000 0.085000 0.310000 0.255000 ;
        RECT 0.620000 0.085000 0.690000 0.255000 ;
        RECT 1.030000 0.085000 1.100000 0.320000 ;
        RECT 1.780000 0.085000 1.850000 0.320000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.920000 0.115000 1.240000 ;
      RECT 0.045000 0.850000 0.780000 0.920000 ;
      RECT 0.710000 0.375000 0.780000 0.850000 ;
      RECT 0.045000 0.185000 0.115000 0.850000 ;
      RECT 0.820000 0.975000 0.920000 1.250000 ;
      RECT 0.850000 0.460000 0.920000 0.975000 ;
      RECT 0.850000 0.390000 1.475000 0.460000 ;
      RECT 1.405000 0.460000 1.475000 0.670000 ;
      RECT 0.850000 0.310000 0.920000 0.390000 ;
      RECT 0.820000 0.175000 0.920000 0.310000 ;
      RECT 1.400000 0.875000 1.470000 1.200000 ;
      RECT 1.400000 0.850000 1.910000 0.875000 ;
      RECT 0.985000 0.780000 1.910000 0.850000 ;
      RECT 1.545000 0.740000 1.910000 0.780000 ;
      RECT 0.985000 0.525000 1.055000 0.780000 ;
      RECT 1.545000 0.320000 1.615000 0.740000 ;
      RECT 1.410000 0.185000 1.615000 0.320000 ;
      RECT 1.975000 0.630000 2.045000 1.215000 ;
      RECT 1.705000 0.495000 2.045000 0.630000 ;
      RECT 1.975000 0.185000 2.045000 0.495000 ;
  END
END DLH_X2

MACRO AND2_X1
  CLASS CORE ;
  FOREIGN AND2_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.610000 0.190000 0.700000 1.250000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0954 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.299 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.415000 0.085000 0.485000 0.325000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.910000 0.305000 1.250000 ;
      RECT 0.235000 0.840000 0.540000 0.910000 ;
      RECT 0.470000 0.460000 0.540000 0.840000 ;
      RECT 0.045000 0.390000 0.540000 0.460000 ;
      RECT 0.045000 0.190000 0.115000 0.390000 ;
  END
END AND2_X1

MACRO AND2_X2
  CLASS CORE ;
  FOREIGN AND2_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.380000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.615000 0.150000 0.700000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.910000 0.305000 1.250000 ;
      RECT 0.235000 0.840000 0.545000 0.910000 ;
      RECT 0.475000 0.460000 0.545000 0.840000 ;
      RECT 0.045000 0.390000 0.545000 0.460000 ;
      RECT 0.045000 0.150000 0.115000 0.390000 ;
  END
END AND2_X2

MACRO AND2_X4
  CLASS CORE ;
  FOREIGN AND2_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.420000 0.380000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0312 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0962 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.420000 0.185000 0.725000 ;
        RECT 0.060000 0.725000 0.760000 0.795000 ;
        RECT 0.690000 0.525000 0.760000 0.725000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.101125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3315 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.150000 1.080000 0.680000 ;
        RECT 0.995000 0.680000 1.435000 0.750000 ;
        RECT 0.995000 0.750000 1.080000 1.250000 ;
        RECT 1.365000 0.750000 1.435000 1.250000 ;
        RECT 1.365000 0.150000 1.435000 0.680000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.19045 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6682 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.040000 0.995000 0.110000 1.315000 ;
        RECT 0.415000 0.995000 0.485000 1.315000 ;
        RECT 0.795000 0.995000 0.865000 1.315000 ;
        RECT 1.175000 0.995000 1.245000 1.315000 ;
        RECT 1.555000 0.995000 1.625000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.355000 ;
        RECT 0.795000 0.085000 0.865000 0.215000 ;
        RECT 1.175000 0.085000 1.245000 0.355000 ;
        RECT 1.555000 0.085000 1.625000 0.355000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.930000 0.305000 1.250000 ;
      RECT 0.235000 0.860000 0.920000 0.930000 ;
      RECT 0.605000 0.930000 0.675000 1.250000 ;
      RECT 0.850000 0.355000 0.920000 0.860000 ;
      RECT 0.425000 0.285000 0.920000 0.355000 ;
      RECT 0.425000 0.220000 0.495000 0.285000 ;
  END
END AND2_X4

MACRO AND3_X1
  CLASS CORE ;
  FOREIGN AND3_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.570000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.800000 0.975000 0.890000 1.250000 ;
        RECT 0.820000 0.425000 0.890000 0.975000 ;
        RECT 0.800000 0.150000 0.890000 0.425000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.088 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3146 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.225000 1.040000 0.295000 1.315000 ;
        RECT 0.605000 1.000000 0.675000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.935000 0.115000 1.250000 ;
      RECT 0.045000 0.865000 0.705000 0.935000 ;
      RECT 0.415000 0.935000 0.485000 1.250000 ;
      RECT 0.635000 0.660000 0.705000 0.865000 ;
      RECT 0.635000 0.525000 0.755000 0.660000 ;
      RECT 0.635000 0.420000 0.705000 0.525000 ;
      RECT 0.045000 0.350000 0.705000 0.420000 ;
      RECT 0.045000 0.150000 0.115000 0.350000 ;
  END
END AND3_X1

MACRO AND3_X2
  CLASS CORE ;
  FOREIGN AND3_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.570000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.805000 0.150000 0.890000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.225000 0.975000 0.295000 1.315000 ;
        RECT 0.605000 0.975000 0.675000 1.315000 ;
        RECT 0.990000 0.975000 1.060000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.605000 0.085000 0.675000 0.285000 ;
        RECT 0.990000 0.085000 1.060000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.870000 0.115000 1.250000 ;
      RECT 0.045000 0.800000 0.735000 0.870000 ;
      RECT 0.415000 0.870000 0.485000 1.250000 ;
      RECT 0.665000 0.425000 0.735000 0.800000 ;
      RECT 0.045000 0.355000 0.735000 0.425000 ;
      RECT 0.045000 0.150000 0.115000 0.355000 ;
  END
END AND3_X2

MACRO AND3_X4
  CLASS CORE ;
  FOREIGN AND3_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.595000 0.555000 0.730000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.019575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.340000 0.420000 0.950000 0.490000 ;
        RECT 0.340000 0.490000 0.410000 0.660000 ;
        RECT 0.820000 0.490000 0.950000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0819 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2756 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.190000 0.700000 ;
        RECT 0.120000 0.700000 0.190000 0.765000 ;
        RECT 0.120000 0.765000 1.140000 0.835000 ;
        RECT 1.070000 0.525000 1.140000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.1155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4238 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.375000 0.150000 1.445000 0.560000 ;
        RECT 1.375000 0.560000 1.815000 0.700000 ;
        RECT 1.375000 0.700000 1.445000 1.250000 ;
        RECT 1.745000 0.700000 1.815000 1.250000 ;
        RECT 1.745000 0.150000 1.815000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.65 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 0.040000 1.035000 0.110000 1.315000 ;
        RECT 0.415000 1.035000 0.485000 1.315000 ;
        RECT 0.795000 1.035000 0.865000 1.315000 ;
        RECT 1.175000 1.035000 1.245000 1.315000 ;
        RECT 1.555000 1.035000 1.625000 1.315000 ;
        RECT 1.935000 1.035000 2.005000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 1.175000 0.085000 1.245000 0.195000 ;
        RECT 1.555000 0.085000 1.625000 0.425000 ;
        RECT 1.935000 0.085000 2.005000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.970000 0.305000 1.250000 ;
      RECT 0.235000 0.900000 1.305000 0.970000 ;
      RECT 0.605000 0.970000 0.675000 1.250000 ;
      RECT 0.985000 0.970000 1.055000 1.250000 ;
      RECT 1.235000 0.330000 1.305000 0.900000 ;
      RECT 0.615000 0.260000 1.305000 0.330000 ;
      RECT 0.615000 0.150000 0.685000 0.260000 ;
  END
END AND3_X4

MACRO AND4_X1
  CLASS CORE ;
  FOREIGN AND4_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.760000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.990000 0.150000 1.080000 1.250000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.099 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3094 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.795000 0.085000 0.865000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.910000 0.305000 1.250000 ;
      RECT 0.235000 0.840000 0.925000 0.910000 ;
      RECT 0.605000 0.910000 0.675000 1.250000 ;
      RECT 0.855000 0.420000 0.925000 0.840000 ;
      RECT 0.045000 0.350000 0.925000 0.420000 ;
      RECT 0.045000 0.150000 0.115000 0.350000 ;
  END
END AND4_X1

MACRO AND4_X2
  CLASS CORE ;
  FOREIGN AND4_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.760000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.150000 1.080000 1.250000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.0935 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3081 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.040000 0.975000 0.110000 1.315000 ;
        RECT 0.415000 0.975000 0.485000 1.315000 ;
        RECT 0.795000 0.975000 0.865000 1.315000 ;
        RECT 1.180000 0.975000 1.250000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.795000 0.085000 0.865000 0.270000 ;
        RECT 1.180000 0.085000 1.250000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.870000 0.305000 1.250000 ;
      RECT 0.235000 0.800000 0.925000 0.870000 ;
      RECT 0.605000 0.870000 0.675000 1.250000 ;
      RECT 0.855000 0.425000 0.925000 0.800000 ;
      RECT 0.045000 0.355000 0.925000 0.425000 ;
      RECT 0.045000 0.150000 0.115000 0.355000 ;
  END
END AND4_X2

MACRO AND4_X4
  CLASS CORE ;
  FOREIGN AND4_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.800000 0.560000 0.935000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.565000 0.425000 1.135000 0.495000 ;
        RECT 0.565000 0.495000 0.700000 0.700000 ;
        RECT 1.065000 0.495000 1.135000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.079125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2626 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.355000 0.525000 0.425000 0.770000 ;
        RECT 0.355000 0.770000 1.345000 0.840000 ;
        RECT 1.200000 0.525000 1.345000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.121975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.403 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A3

  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.205000 0.700000 ;
        RECT 0.135000 0.700000 0.205000 0.905000 ;
        RECT 0.135000 0.905000 1.535000 0.975000 ;
        RECT 1.465000 0.525000 1.535000 0.905000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.164325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5993 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A4

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.770000 0.150000 1.840000 0.560000 ;
        RECT 1.770000 0.560000 2.210000 0.700000 ;
        RECT 1.770000 0.700000 1.840000 0.925000 ;
        RECT 2.140000 0.700000 2.210000 0.925000 ;
        RECT 2.140000 0.150000 2.210000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1505 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.481 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.430000 1.175000 0.500000 1.315000 ;
        RECT 0.810000 1.175000 0.880000 1.315000 ;
        RECT 1.190000 1.175000 1.260000 1.315000 ;
        RECT 1.570000 1.175000 1.640000 1.315000 ;
        RECT 0.055000 1.065000 0.125000 1.315000 ;
        RECT 1.950000 1.065000 2.020000 1.315000 ;
        RECT 2.330000 1.065000 2.400000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.425000 ;
        RECT 1.570000 0.085000 1.640000 0.195000 ;
        RECT 1.950000 0.085000 2.020000 0.425000 ;
        RECT 2.330000 0.085000 2.400000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215000 1.040000 1.705000 1.110000 ;
      RECT 1.635000 0.360000 1.705000 1.040000 ;
      RECT 0.785000 0.290000 1.705000 0.360000 ;
  END
END AND4_X4

MACRO ANTENNA_X1
  CLASS CORE ;
  FOREIGN ANTENNA_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.19 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.420000 0.130000 0.750000 ;
    END
    ANTENNAGATEAREA 0.0162 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0231 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.104 LAYER metal1 ;
    ANTENNAGATEAREA 0.0162 LAYER metal2 ;
    ANTENNAGATEAREA 0.0162 LAYER metal3 ;
    ANTENNAGATEAREA 0.0162 LAYER metal4 ;
    ANTENNAGATEAREA 0.0162 LAYER metal5 ;
    ANTENNAGATEAREA 0.0162 LAYER metal6 ;
    ANTENNAGATEAREA 0.0162 LAYER metal7 ;
    ANTENNAGATEAREA 0.0162 LAYER metal8 ;
    ANTENNAGATEAREA 0.0162 LAYER metal9 ;
    ANTENNAGATEAREA 0.0162 LAYER metal10 ;
  END A

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.190000 1.485000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.190000 0.085000 ;
    END
  END VSS
END ANTENNA_X1

MACRO AOI211_X1
  CLASS CORE ;
  FOREIGN AOI211_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.410000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.210000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0845 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.275000 0.355000 0.905000 0.425000 ;
        RECT 0.275000 0.425000 0.345000 1.115000 ;
        RECT 0.440000 0.150000 0.525000 0.355000 ;
        RECT 0.835000 0.150000 0.905000 0.355000 ;
    END
    ANTENNADIFFAREA 0.189875 ;
    ANTENNAPARTIALMETALAREA 0.124175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.468 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.835000 0.905000 0.905000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.425000 ;
        RECT 0.645000 0.085000 0.715000 0.285000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085000 1.180000 0.525000 1.250000 ;
      RECT 0.085000 0.905000 0.155000 1.180000 ;
      RECT 0.455000 0.905000 0.525000 1.180000 ;
  END
END AOI211_X1

MACRO AOI211_X2
  CLASS CORE ;
  FOREIGN AOI211_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.390000 0.560000 0.525000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.765000 ;
        RECT 0.060000 0.765000 0.750000 0.835000 ;
        RECT 0.680000 0.525000 0.750000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0951 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3224 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.190000 0.560000 1.325000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.965000 0.425000 1.650000 0.495000 ;
        RECT 0.965000 0.495000 1.035000 0.660000 ;
        RECT 1.540000 0.495000 1.650000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08205 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2925 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.355000 0.890000 0.765000 ;
        RECT 0.820000 0.765000 1.475000 0.835000 ;
        RECT 0.200000 0.285000 1.320000 0.355000 ;
        RECT 1.025000 0.835000 1.095000 1.055000 ;
        RECT 1.405000 0.835000 1.475000 1.055000 ;
        RECT 0.200000 0.150000 0.335000 0.285000 ;
        RECT 1.185000 0.150000 1.320000 0.285000 ;
    END
    ANTENNADIFFAREA 0.3507 ;
    ANTENNAPARTIALMETALAREA 0.2202 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7709 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.420000 1.035000 0.490000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.045000 0.085000 0.115000 0.355000 ;
        RECT 0.430000 0.085000 0.500000 0.215000 ;
        RECT 0.825000 0.085000 0.895000 0.215000 ;
        RECT 1.595000 0.085000 1.665000 0.355000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.815000 1.180000 1.665000 1.250000 ;
      RECT 1.220000 0.975000 1.290000 1.180000 ;
      RECT 1.595000 0.975000 1.665000 1.180000 ;
      RECT 0.815000 0.970000 0.885000 1.180000 ;
      RECT 0.050000 0.900000 0.885000 0.970000 ;
      RECT 0.050000 0.970000 0.120000 1.250000 ;
  END
END AOI211_X2

MACRO AOI211_X4
  CLASS CORE ;
  FOREIGN AOI211_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.760000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.375000 0.150000 1.445000 0.560000 ;
        RECT 1.375000 0.560000 1.820000 0.700000 ;
        RECT 1.375000 0.700000 1.445000 1.175000 ;
        RECT 1.750000 0.700000 1.820000 1.175000 ;
        RECT 1.750000 0.150000 1.820000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.1862 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6123 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 0.795000 0.900000 0.865000 1.315000 ;
        RECT 1.175000 0.900000 1.245000 1.315000 ;
        RECT 1.555000 0.900000 1.625000 1.315000 ;
        RECT 1.935000 0.900000 2.005000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.415000 0.085000 0.485000 0.285000 ;
        RECT 0.795000 0.085000 0.865000 0.285000 ;
        RECT 1.175000 0.085000 1.245000 0.425000 ;
        RECT 1.555000 0.085000 1.625000 0.425000 ;
        RECT 1.935000 0.085000 2.005000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 1.180000 0.485000 1.250000 ;
      RECT 0.045000 0.900000 0.115000 1.180000 ;
      RECT 0.415000 0.900000 0.485000 1.180000 ;
      RECT 0.235000 0.835000 0.305000 1.115000 ;
      RECT 0.235000 0.765000 0.930000 0.835000 ;
      RECT 0.860000 0.460000 0.930000 0.765000 ;
      RECT 0.045000 0.390000 0.930000 0.460000 ;
      RECT 0.045000 0.150000 0.115000 0.390000 ;
      RECT 0.605000 0.150000 0.675000 0.390000 ;
      RECT 0.995000 0.660000 1.065000 1.175000 ;
      RECT 0.995000 0.525000 1.310000 0.660000 ;
      RECT 0.995000 0.150000 1.065000 0.525000 ;
  END
END AOI211_X4

MACRO AOI21_X1
  CLASS CORE ;
  FOREIGN AOI21_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.76 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.400000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.200000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0819 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.265000 0.355000 0.525000 0.425000 ;
        RECT 0.265000 0.425000 0.335000 1.115000 ;
        RECT 0.440000 0.150000 0.525000 0.355000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.083925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3185 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.760000 1.485000 ;
        RECT 0.645000 0.905000 0.715000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.760000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.425000 ;
        RECT 0.645000 0.085000 0.715000 0.355000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085000 1.180000 0.525000 1.250000 ;
      RECT 0.085000 0.905000 0.155000 1.180000 ;
      RECT 0.455000 0.905000 0.525000 1.180000 ;
  END
END AOI21_X1

MACRO AOI21_X2
  CLASS CORE ;
  FOREIGN AOI21_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.33 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.215000 0.560000 0.350000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.560000 0.900000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.570000 0.525000 0.700000 0.700000 ;
        RECT 0.630000 0.700000 0.700000 0.770000 ;
        RECT 0.630000 0.770000 1.180000 0.840000 ;
        RECT 1.110000 0.525000 1.180000 0.770000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0833 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3042 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.435000 0.425000 0.505000 0.905000 ;
        RECT 0.435000 0.905000 1.130000 0.975000 ;
        RECT 0.250000 0.355000 0.905000 0.425000 ;
        RECT 0.250000 0.150000 0.335000 0.355000 ;
        RECT 0.835000 0.150000 0.905000 0.355000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.159875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6006 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.330000 1.485000 ;
        RECT 0.265000 1.205000 0.335000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.330000 0.085000 ;
        RECT 0.080000 0.085000 0.150000 0.425000 ;
        RECT 0.455000 0.085000 0.525000 0.285000 ;
        RECT 1.215000 0.085000 1.285000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.085000 1.140000 0.155000 1.250000 ;
      RECT 0.085000 1.070000 1.285000 1.140000 ;
      RECT 1.215000 1.140000 1.285000 1.250000 ;
      RECT 0.085000 0.975000 0.155000 1.070000 ;
      RECT 1.215000 0.975000 1.285000 1.070000 ;
  END
END AOI21_X2

MACRO AOI21_X4
  CLASS CORE ;
  FOREIGN AOI21_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.400000 0.525000 0.535000 0.700000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.023625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.165000 0.560000 1.300000 0.690000 ;
        RECT 1.165000 0.690000 2.060000 0.760000 ;
        RECT 1.925000 0.560000 2.060000 0.690000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09775 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3185 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.925000 0.420000 2.320000 0.490000 ;
        RECT 0.925000 0.490000 0.995000 0.660000 ;
        RECT 1.525000 0.490000 1.660000 0.625000 ;
        RECT 2.250000 0.490000 2.320000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.139675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5044 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.825000 2.210000 0.895000 ;
        RECT 0.630000 0.425000 0.700000 0.825000 ;
        RECT 1.000000 0.895000 1.070000 1.115000 ;
        RECT 1.380000 0.895000 1.450000 1.115000 ;
        RECT 1.760000 0.895000 1.830000 1.115000 ;
        RECT 2.140000 0.895000 2.210000 1.115000 ;
        RECT 0.250000 0.355000 0.700000 0.425000 ;
        RECT 0.630000 0.330000 0.700000 0.355000 ;
        RECT 0.250000 0.150000 0.320000 0.355000 ;
        RECT 0.630000 0.260000 2.055000 0.330000 ;
        RECT 0.630000 0.150000 0.700000 0.260000 ;
    END
    ANTENNADIFFAREA 0.5852 ;
    ANTENNAPARTIALMETALAREA 0.35525 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3377 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.240000 1.205000 0.310000 1.315000 ;
        RECT 0.620000 1.205000 0.690000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.425000 ;
        RECT 0.430000 0.085000 0.500000 0.195000 ;
        RECT 0.810000 0.085000 0.880000 0.195000 ;
        RECT 1.570000 0.085000 1.640000 0.195000 ;
        RECT 2.330000 0.085000 2.400000 0.350000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 1.035000 0.130000 1.240000 ;
      RECT 0.060000 0.965000 0.880000 1.035000 ;
      RECT 0.430000 1.035000 0.500000 1.240000 ;
      RECT 0.810000 1.035000 0.880000 1.180000 ;
      RECT 0.810000 1.180000 2.400000 1.250000 ;
      RECT 1.190000 0.960000 1.260000 1.180000 ;
      RECT 1.570000 0.960000 1.640000 1.180000 ;
      RECT 1.950000 0.960000 2.020000 1.180000 ;
      RECT 2.330000 0.840000 2.400000 1.180000 ;
  END
END AOI21_X4

MACRO AOI221_X1
  CLASS CORE ;
  FOREIGN AOI221_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.14 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.525000 0.565000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.630000 0.525000 0.740000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01925 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0741 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.425000 0.150000 0.495000 0.355000 ;
        RECT 0.425000 0.355000 1.055000 0.425000 ;
        RECT 0.805000 0.425000 0.890000 1.115000 ;
        RECT 0.985000 0.150000 1.055000 0.355000 ;
    END
    ANTENNADIFFAREA 0.189875 ;
    ANTENNAPARTIALMETALAREA 0.13145 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.468 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.140000 1.485000 ;
        RECT 0.225000 0.905000 0.295000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.140000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.355000 ;
        RECT 0.605000 0.085000 0.675000 0.215000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.840000 0.115000 1.180000 ;
      RECT 0.045000 0.770000 0.485000 0.840000 ;
      RECT 0.415000 0.840000 0.485000 1.180000 ;
      RECT 0.615000 1.180000 1.055000 1.250000 ;
      RECT 0.615000 0.905000 0.685000 1.180000 ;
      RECT 0.985000 0.905000 1.055000 1.180000 ;
  END
END AOI221_X1

MACRO AOI221_X2
  CLASS CORE ;
  FOREIGN AOI221_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.09 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.560000 0.250000 0.700000 ;
        RECT 0.180000 0.700000 0.250000 0.790000 ;
        RECT 0.180000 0.790000 1.130000 0.860000 ;
        RECT 1.060000 0.525000 1.130000 0.790000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.11795 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4251 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.340000 0.420000 0.945000 0.490000 ;
        RECT 0.340000 0.490000 0.410000 0.660000 ;
        RECT 0.820000 0.490000 0.945000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0805 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2743 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.585000 0.560000 0.725000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0196 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0728 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.570000 0.525000 1.660000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.340000 0.525000 1.410000 0.765000 ;
        RECT 1.340000 0.765000 1.840000 0.835000 ;
        RECT 1.770000 0.700000 1.840000 0.765000 ;
        RECT 1.770000 0.525000 1.910000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08085 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2912 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.195000 0.900000 1.860000 0.970000 ;
        RECT 1.195000 0.350000 1.275000 0.900000 ;
        RECT 0.200000 0.280000 1.675000 0.350000 ;
    END
    ANTENNADIFFAREA 0.3507 ;
    ANTENNAPARTIALMETALAREA 0.1938 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.715 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.090000 1.485000 ;
        RECT 0.415000 1.205000 0.485000 1.315000 ;
        RECT 0.795000 1.205000 0.865000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.090000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.425000 ;
        RECT 0.605000 0.085000 0.675000 0.195000 ;
        RECT 1.175000 0.085000 1.245000 0.195000 ;
        RECT 1.945000 0.085000 2.015000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200000 0.930000 1.090000 1.000000 ;
      RECT 0.045000 1.070000 2.015000 1.140000 ;
      RECT 0.045000 0.865000 0.115000 1.070000 ;
      RECT 1.945000 0.865000 2.015000 1.070000 ;
  END
END AOI221_X2

MACRO AOI221_X4
  CLASS CORE ;
  FOREIGN AOI221_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.47 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.610000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.800000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.180000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02975 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0897 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.270000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.03675 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1001 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.420000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.795000 0.150000 1.885000 0.560000 ;
        RECT 1.795000 0.560000 2.240000 0.700000 ;
        RECT 1.795000 0.700000 1.865000 1.250000 ;
        RECT 2.170000 0.700000 2.240000 1.250000 ;
        RECT 2.170000 0.150000 2.240000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.2049 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6513 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.470000 1.485000 ;
        RECT 0.875000 1.035000 0.945000 1.315000 ;
        RECT 1.600000 1.005000 1.670000 1.315000 ;
        RECT 1.215000 0.975000 1.285000 1.315000 ;
        RECT 1.975000 0.975000 2.045000 1.315000 ;
        RECT 2.355000 0.975000 2.425000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.470000 0.085000 ;
        RECT 0.495000 0.085000 0.565000 0.285000 ;
        RECT 1.215000 0.085000 1.285000 0.285000 ;
        RECT 1.605000 0.085000 1.675000 0.425000 ;
        RECT 1.975000 0.085000 2.045000 0.425000 ;
        RECT 2.355000 0.085000 2.425000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.125000 1.175000 0.195000 1.250000 ;
      RECT 0.125000 1.105000 0.565000 1.175000 ;
      RECT 0.495000 1.175000 0.565000 1.250000 ;
      RECT 0.125000 0.975000 0.195000 1.105000 ;
      RECT 0.495000 0.975000 0.565000 1.105000 ;
      RECT 0.695000 0.970000 0.765000 1.250000 ;
      RECT 0.695000 0.900000 1.100000 0.970000 ;
      RECT 1.030000 0.970000 1.100000 1.250000 ;
      RECT 0.315000 0.835000 0.385000 1.040000 ;
      RECT 0.315000 0.765000 1.350000 0.835000 ;
      RECT 1.280000 0.425000 1.350000 0.765000 ;
      RECT 0.125000 0.355000 1.350000 0.425000 ;
      RECT 0.125000 0.150000 0.195000 0.355000 ;
      RECT 0.710000 0.150000 0.780000 0.355000 ;
      RECT 1.415000 0.660000 1.485000 1.250000 ;
      RECT 1.415000 0.525000 1.730000 0.660000 ;
      RECT 1.415000 0.150000 1.485000 0.525000 ;
  END
END AOI221_X4

MACRO AOI222_X1
  CLASS CORE ;
  FOREIGN AOI222_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.52 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.315000 0.525000 1.460000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.025375 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0832 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.995000 0.525000 1.080000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.014875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0676 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.620000 0.525000 0.720000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.525000 0.910000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.01575 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0689 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.215000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.027125 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0858 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.500000 0.175000 0.570000 0.375000 ;
        RECT 0.500000 0.375000 1.460000 0.450000 ;
        RECT 1.145000 0.450000 1.215000 1.115000 ;
        RECT 1.325000 0.175000 1.460000 0.375000 ;
    END
    ANTENNADIFFAREA 0.252125 ;
    ANTENNAPARTIALMETALAREA 0.15955 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.546 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.520000 1.485000 ;
        RECT 0.040000 0.905000 0.110000 1.315000 ;
        RECT 0.415000 0.905000 0.485000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.520000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.450000 ;
        RECT 0.945000 0.085000 1.015000 0.310000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235000 0.840000 0.305000 1.180000 ;
      RECT 0.235000 0.770000 0.825000 0.840000 ;
      RECT 0.755000 0.840000 0.825000 1.115000 ;
      RECT 0.575000 1.180000 1.395000 1.250000 ;
      RECT 0.575000 0.905000 0.645000 1.180000 ;
      RECT 0.945000 0.905000 1.015000 1.180000 ;
      RECT 1.325000 0.905000 1.395000 1.180000 ;
  END
END AOI222_X1

MACRO AOI222_X2
  CLASS CORE ;
  FOREIGN AOI222_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.910000 0.560000 2.045000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 2.285000 0.560000 2.420000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.145000 0.560000 1.280000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.910000 0.420000 1.545000 0.490000 ;
        RECT 0.910000 0.490000 1.080000 0.660000 ;
        RECT 1.475000 0.490000 1.545000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.08525 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2717 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.560000 0.520000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.425000 0.760000 0.495000 ;
        RECT 0.060000 0.495000 0.190000 0.700000 ;
        RECT 0.690000 0.495000 0.760000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0872 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2964 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.770000 0.770000 2.380000 0.840000 ;
        RECT 1.770000 0.355000 1.840000 0.770000 ;
        RECT 1.940000 0.840000 2.010000 1.115000 ;
        RECT 2.310000 0.840000 2.380000 1.115000 ;
        RECT 0.390000 0.285000 2.035000 0.355000 ;
        RECT 0.390000 0.150000 0.525000 0.285000 ;
        RECT 1.145000 0.150000 1.280000 0.285000 ;
    END
    ANTENNADIFFAREA 0.3507 ;
    ANTENNAPARTIALMETALAREA 0.26185 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.9256 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.660000 1.485000 ;
        RECT 0.225000 0.905000 0.295000 1.315000 ;
        RECT 0.605000 0.905000 0.675000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.660000 0.085000 ;
        RECT 0.040000 0.085000 0.110000 0.250000 ;
        RECT 0.765000 0.085000 0.900000 0.215000 ;
        RECT 1.555000 0.085000 1.625000 0.195000 ;
        RECT 2.310000 0.085000 2.380000 0.250000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.840000 0.115000 1.180000 ;
      RECT 0.045000 0.770000 1.625000 0.840000 ;
      RECT 0.415000 0.840000 0.485000 1.180000 ;
      RECT 0.795000 0.840000 0.865000 1.180000 ;
      RECT 1.175000 0.840000 1.245000 1.115000 ;
      RECT 1.555000 0.840000 1.625000 1.115000 ;
      RECT 2.100000 0.355000 2.570000 0.425000 ;
      RECT 2.100000 0.220000 2.170000 0.355000 ;
      RECT 2.500000 0.150000 2.570000 0.355000 ;
      RECT 1.715000 0.150000 2.170000 0.220000 ;
      RECT 0.995000 1.180000 2.570000 1.250000 ;
      RECT 0.995000 0.905000 1.065000 1.180000 ;
      RECT 1.365000 0.905000 1.435000 1.180000 ;
      RECT 1.745000 0.905000 1.815000 1.180000 ;
      RECT 2.120000 0.905000 2.190000 1.180000 ;
      RECT 2.500000 0.905000 2.570000 1.180000 ;
  END
END AOI222_X2

MACRO AOI222_X4
  CLASS CORE ;
  FOREIGN AOI222_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 2.66 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.235000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.030625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.091 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.385000 0.525000 0.510000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.525000 0.890000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.525000 0.700000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.010000 0.525000 1.135000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C1

  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.200000 0.525000 1.335000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.023625 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0806 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END C2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.950000 0.150000 2.020000 0.560000 ;
        RECT 1.950000 0.560000 2.410000 0.700000 ;
        RECT 1.950000 0.700000 2.020000 1.205000 ;
        RECT 2.330000 0.700000 2.410000 1.205000 ;
        RECT 2.325000 0.150000 2.410000 0.560000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.2037 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6318 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 2.660000 1.485000 ;
        RECT 0.995000 1.065000 1.065000 1.315000 ;
        RECT 1.370000 0.930000 1.440000 1.315000 ;
        RECT 1.750000 0.930000 1.820000 1.315000 ;
        RECT 2.130000 0.930000 2.200000 1.315000 ;
        RECT 2.510000 0.930000 2.580000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 2.660000 0.085000 ;
        RECT 0.460000 0.085000 0.530000 0.285000 ;
        RECT 1.370000 0.085000 1.440000 0.285000 ;
        RECT 1.750000 0.085000 1.820000 0.425000 ;
        RECT 2.140000 0.085000 2.210000 0.425000 ;
        RECT 2.510000 0.085000 2.580000 0.425000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.090000 1.135000 0.910000 1.205000 ;
      RECT 0.840000 1.070000 0.910000 1.135000 ;
      RECT 0.090000 0.930000 0.160000 1.135000 ;
      RECT 0.460000 0.930000 0.530000 1.135000 ;
      RECT 0.660000 1.000000 0.730000 1.065000 ;
      RECT 0.660000 0.930000 1.250000 1.000000 ;
      RECT 1.180000 1.000000 1.250000 1.205000 ;
      RECT 0.280000 0.835000 0.350000 1.040000 ;
      RECT 0.280000 0.765000 1.505000 0.835000 ;
      RECT 1.435000 0.425000 1.505000 0.765000 ;
      RECT 0.090000 0.355000 1.505000 0.425000 ;
      RECT 0.090000 0.150000 0.160000 0.355000 ;
      RECT 0.840000 0.150000 0.910000 0.355000 ;
      RECT 1.570000 0.660000 1.640000 1.205000 ;
      RECT 1.570000 0.525000 1.885000 0.660000 ;
      RECT 1.570000 0.150000 1.640000 0.525000 ;
  END
END AOI222_X4

MACRO AOI22_X1
  CLASS CORE ;
  FOREIGN AOI22_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.95 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.575000 0.420000 0.700000 0.660000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.03 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0949 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.765000 0.420000 0.890000 0.660000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.03 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0949 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.250000 0.525000 0.375000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.185000 0.700000 ;
    END
    ANTENNAGATEAREA 0.05225 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.021875 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.078 LAYER metal1 ;
    ANTENNAGATEAREA 0.05225 LAYER metal2 ;
    ANTENNAGATEAREA 0.05225 LAYER metal3 ;
    ANTENNAGATEAREA 0.05225 LAYER metal4 ;
    ANTENNAGATEAREA 0.05225 LAYER metal5 ;
    ANTENNAGATEAREA 0.05225 LAYER metal6 ;
    ANTENNAGATEAREA 0.05225 LAYER metal7 ;
    ANTENNAGATEAREA 0.05225 LAYER metal8 ;
    ANTENNAGATEAREA 0.05225 LAYER metal9 ;
    ANTENNAGATEAREA 0.05225 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.440000 0.150000 0.510000 0.725000 ;
        RECT 0.440000 0.725000 0.690000 0.795000 ;
        RECT 0.620000 0.795000 0.690000 1.005000 ;
    END
    ANTENNADIFFAREA 0.1463 ;
    ANTENNAPARTIALMETALAREA 0.07245 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2873 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.950000 1.485000 ;
        RECT 0.240000 1.205000 0.310000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.950000 0.085000 ;
        RECT 0.055000 0.085000 0.125000 0.355000 ;
        RECT 0.810000 0.085000 0.880000 0.355000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.060000 1.070000 0.880000 1.140000 ;
      RECT 0.060000 0.865000 0.130000 1.070000 ;
      RECT 0.435000 0.865000 0.505000 1.070000 ;
      RECT 0.810000 0.865000 0.880000 1.070000 ;
  END
END AOI22_X1

MACRO AOI22_X2
  CLASS CORE ;
  FOREIGN AOI22_X2 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 1.71 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.155000 0.560000 1.290000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.955000 0.425000 1.550000 0.495000 ;
        RECT 0.955000 0.495000 1.080000 0.700000 ;
        RECT 1.480000 0.495000 1.550000 0.660000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.078825 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2691 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395000 0.560000 0.530000 0.700000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.0189 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0715 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.195000 0.765000 ;
        RECT 0.060000 0.765000 0.755000 0.835000 ;
        RECT 0.685000 0.525000 0.755000 0.765000 ;
    END
    ANTENNAGATEAREA 0.1045 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09785 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3237 LAYER metal1 ;
    ANTENNAGATEAREA 0.1045 LAYER metal2 ;
    ANTENNAGATEAREA 0.1045 LAYER metal3 ;
    ANTENNAGATEAREA 0.1045 LAYER metal4 ;
    ANTENNAGATEAREA 0.1045 LAYER metal5 ;
    ANTENNAGATEAREA 0.1045 LAYER metal6 ;
    ANTENNAGATEAREA 0.1045 LAYER metal7 ;
    ANTENNAGATEAREA 0.1045 LAYER metal8 ;
    ANTENNAGATEAREA 0.1045 LAYER metal9 ;
    ANTENNAGATEAREA 0.1045 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.820000 0.355000 0.890000 0.765000 ;
        RECT 0.820000 0.765000 1.445000 0.835000 ;
        RECT 0.395000 0.280000 1.285000 0.355000 ;
        RECT 0.990000 0.835000 1.060000 1.065000 ;
        RECT 1.375000 0.835000 1.445000 1.065000 ;
        RECT 0.395000 0.150000 0.530000 0.280000 ;
        RECT 1.150000 0.150000 1.285000 0.280000 ;
    END
    ANTENNADIFFAREA 0.2926 ;
    ANTENNAPARTIALMETALAREA 0.2065 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7072 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 1.710000 1.485000 ;
        RECT 0.230000 1.035000 0.300000 1.315000 ;
        RECT 0.610000 1.035000 0.680000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 1.710000 0.085000 ;
        RECT 0.045000 0.085000 0.115000 0.390000 ;
        RECT 0.770000 0.085000 0.905000 0.205000 ;
        RECT 1.560000 0.085000 1.630000 0.360000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.800000 1.180000 1.630000 1.250000 ;
      RECT 1.180000 0.975000 1.250000 1.180000 ;
      RECT 1.560000 0.975000 1.630000 1.180000 ;
      RECT 0.800000 0.970000 0.870000 1.180000 ;
      RECT 0.050000 0.900000 0.870000 0.970000 ;
      RECT 0.050000 0.970000 0.120000 1.250000 ;
      RECT 0.420000 0.970000 0.490000 1.250000 ;
  END
END AOI22_X2

MACRO AOI22_X4
  CLASS CORE ;
  FOREIGN AOI22_X4 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 3.23 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.915000 0.560000 2.050000 0.690000 ;
        RECT 1.915000 0.690000 2.790000 0.760000 ;
        RECT 2.655000 0.560000 2.790000 0.690000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09635 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3133 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A1

  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.715000 0.420000 3.045000 0.490000 ;
        RECT 1.715000 0.490000 1.785000 0.660000 ;
        RECT 2.295000 0.490000 2.430000 0.625000 ;
        RECT 2.910000 0.490000 3.045000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.146175 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4875 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END A2

  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.395000 0.560000 0.530000 0.690000 ;
        RECT 0.395000 0.690000 1.290000 0.760000 ;
        RECT 1.155000 0.560000 1.290000 0.690000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.09775 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3185 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B1

  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.125000 0.420000 1.515000 0.490000 ;
        RECT 0.125000 0.490000 0.195000 0.660000 ;
        RECT 0.755000 0.490000 0.890000 0.625000 ;
        RECT 1.445000 0.490000 1.515000 0.660000 ;
    END
    ANTENNAGATEAREA 0.209 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.139325 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.5031 LAYER metal1 ;
    ANTENNAGATEAREA 0.209 LAYER metal2 ;
    ANTENNAGATEAREA 0.209 LAYER metal3 ;
    ANTENNAGATEAREA 0.209 LAYER metal4 ;
    ANTENNAGATEAREA 0.209 LAYER metal5 ;
    ANTENNAGATEAREA 0.209 LAYER metal6 ;
    ANTENNAGATEAREA 0.209 LAYER metal7 ;
    ANTENNAGATEAREA 0.209 LAYER metal8 ;
    ANTENNAGATEAREA 0.209 LAYER metal9 ;
    ANTENNAGATEAREA 0.209 LAYER metal10 ;
  END B2

  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.580000 0.725000 1.820000 0.795000 ;
        RECT 1.580000 0.330000 1.650000 0.725000 ;
        RECT 1.750000 0.795000 1.820000 0.825000 ;
        RECT 0.395000 0.260000 2.805000 0.330000 ;
        RECT 1.750000 0.825000 2.960000 0.895000 ;
        RECT 1.750000 0.895000 1.820000 1.115000 ;
        RECT 2.130000 0.895000 2.200000 1.115000 ;
        RECT 2.510000 0.895000 2.580000 1.115000 ;
        RECT 2.890000 0.895000 2.960000 1.115000 ;
    END
    ANTENNADIFFAREA 0.5852 ;
    ANTENNAPARTIALMETALAREA 0.36155 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3611 LAYER metal1 ;
  END ZN

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 3.230000 1.485000 ;
        RECT 0.230000 1.065000 0.300000 1.315000 ;
        RECT 0.610000 1.065000 0.680000 1.315000 ;
        RECT 0.990000 1.065000 1.060000 1.315000 ;
        RECT 1.370000 1.065000 1.440000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 3.230000 0.085000 ;
        RECT 0.045000 0.085000 0.115000 0.335000 ;
        RECT 0.770000 0.085000 0.905000 0.160000 ;
        RECT 1.530000 0.085000 1.665000 0.160000 ;
        RECT 2.290000 0.085000 2.425000 0.160000 ;
        RECT 3.080000 0.085000 3.150000 0.335000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 1.560000 1.180000 3.150000 1.250000 ;
      RECT 1.940000 0.960000 2.010000 1.180000 ;
      RECT 2.320000 0.960000 2.390000 1.180000 ;
      RECT 2.700000 0.960000 2.770000 1.180000 ;
      RECT 1.560000 0.940000 1.630000 1.180000 ;
      RECT 3.080000 0.840000 3.150000 1.180000 ;
      RECT 0.050000 0.870000 1.630000 0.940000 ;
      RECT 0.050000 0.940000 0.120000 1.160000 ;
      RECT 0.420000 0.940000 0.490000 1.160000 ;
      RECT 0.800000 0.940000 0.870000 1.160000 ;
      RECT 1.180000 0.940000 1.250000 1.160000 ;
  END
END AOI22_X4

MACRO BUF_X1
  CLASS CORE ;
  FOREIGN BUF_X1 0 0 N ;
  ORIGIN 0 0 ;
  SIZE 0.57 BY 1.4 ;
  SYMMETRY X Y ;
  SITE unit ;

  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.060000 0.525000 0.190000 0.700000 ;
    END
    ANTENNAGATEAREA 0.02625 LAYER metal1 ;
    ANTENNAPARTIALMETALAREA 0.02275 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0793 LAYER metal1 ;
    ANTENNAGATEAREA 0.02625 LAYER metal2 ;
    ANTENNAGATEAREA 0.02625 LAYER metal3 ;
    ANTENNAGATEAREA 0.02625 LAYER metal4 ;
    ANTENNAGATEAREA 0.02625 LAYER metal5 ;
    ANTENNAGATEAREA 0.02625 LAYER metal6 ;
    ANTENNAGATEAREA 0.02625 LAYER metal7 ;
    ANTENNAGATEAREA 0.02625 LAYER metal8 ;
    ANTENNAGATEAREA 0.02625 LAYER metal9 ;
    ANTENNAGATEAREA 0.02625 LAYER metal10 ;
  END A

  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.420000 0.190000 0.510000 1.240000 ;
    END
    ANTENNADIFFAREA 0.109725 ;
    ANTENNAPARTIALMETALAREA 0.0945 LAYER metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2964 LAYER metal1 ;
  END Z

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 1.315000 0.570000 1.485000 ;
        RECT 0.225000 0.965000 0.295000 1.315000 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.000000 -0.085000 0.570000 0.085000 ;
        RECT 0.225000 0.085000 0.295000 0.325000 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045000 0.900000 0.115000 1.240000 ;
      RECT 0.045000 0.830000 0.355000 0.900000 ;
      RECT 0.285000 0.460000 0.355000 0.830000 ;
      RECT 0.045000 0.390000 0.355000 0.460000 ;
      RECT 0.045000 0.190000 0.115000 0.390000 ;
  END
END BUF_X1
  
END LIBRARY
